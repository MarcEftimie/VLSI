magic
tech sky130A
timestamp 1695601967
<< nwell >>
rect 85 -405 470 440
<< nmos >>
rect 250 -540 265 -440
rect 250 -690 265 -590
rect 185 -795 315 -780
rect 185 -860 315 -845
rect 185 -925 315 -910
rect 210 -1070 310 -1055
rect 210 -1135 310 -1120
rect 210 -1280 310 -1265
rect 210 -1345 310 -1330
<< pmos >>
rect 210 350 310 365
rect 210 285 310 300
rect 210 140 310 155
rect 210 75 310 90
rect 250 -105 265 -5
rect 250 -235 265 -135
rect 250 -385 265 -285
<< ndiff >>
rect 200 -455 250 -440
rect 200 -525 215 -455
rect 235 -525 250 -455
rect 200 -540 250 -525
rect 265 -455 315 -440
rect 265 -525 280 -455
rect 300 -525 315 -455
rect 265 -540 315 -525
rect 200 -605 250 -590
rect 200 -675 215 -605
rect 235 -675 250 -605
rect 200 -690 250 -675
rect 265 -605 315 -590
rect 265 -675 280 -605
rect 300 -675 315 -605
rect 265 -690 315 -675
rect 185 -745 315 -730
rect 185 -765 200 -745
rect 300 -765 315 -745
rect 185 -780 315 -765
rect 185 -810 315 -795
rect 185 -830 200 -810
rect 300 -830 315 -810
rect 185 -845 315 -830
rect 185 -875 315 -860
rect 185 -895 200 -875
rect 300 -895 315 -875
rect 185 -910 315 -895
rect 185 -940 315 -925
rect 185 -960 200 -940
rect 300 -960 315 -940
rect 185 -975 315 -960
rect 210 -1020 310 -1005
rect 210 -1040 225 -1020
rect 295 -1040 310 -1020
rect 210 -1055 310 -1040
rect 210 -1085 310 -1070
rect 210 -1105 225 -1085
rect 295 -1105 310 -1085
rect 210 -1120 310 -1105
rect 210 -1150 310 -1135
rect 210 -1170 225 -1150
rect 295 -1170 310 -1150
rect 210 -1185 310 -1170
rect 210 -1230 310 -1215
rect 210 -1250 225 -1230
rect 295 -1250 310 -1230
rect 210 -1265 310 -1250
rect 210 -1295 310 -1280
rect 210 -1315 225 -1295
rect 295 -1315 310 -1295
rect 210 -1330 310 -1315
rect 210 -1360 310 -1345
rect 210 -1380 225 -1360
rect 295 -1380 310 -1360
rect 210 -1395 310 -1380
<< pdiff >>
rect 210 400 310 415
rect 210 380 225 400
rect 295 380 310 400
rect 210 365 310 380
rect 210 335 310 350
rect 210 315 225 335
rect 295 315 310 335
rect 210 300 310 315
rect 210 270 310 285
rect 210 250 225 270
rect 295 250 310 270
rect 210 235 310 250
rect 210 190 310 205
rect 210 170 225 190
rect 295 170 310 190
rect 210 155 310 170
rect 210 125 310 140
rect 210 105 225 125
rect 295 105 310 125
rect 210 90 310 105
rect 210 60 310 75
rect 210 40 225 60
rect 295 40 310 60
rect 210 25 310 40
rect 200 -20 250 -5
rect 200 -90 215 -20
rect 235 -90 250 -20
rect 200 -105 250 -90
rect 265 -20 315 -5
rect 265 -90 280 -20
rect 300 -90 315 -20
rect 265 -105 315 -90
rect 200 -150 250 -135
rect 200 -220 215 -150
rect 235 -220 250 -150
rect 200 -235 250 -220
rect 265 -150 315 -135
rect 265 -220 280 -150
rect 300 -220 315 -150
rect 265 -235 315 -220
rect 200 -300 250 -285
rect 200 -370 215 -300
rect 235 -370 250 -300
rect 200 -385 250 -370
rect 265 -300 315 -285
rect 265 -370 280 -300
rect 300 -370 315 -300
rect 265 -385 315 -370
<< ndiffc >>
rect 215 -525 235 -455
rect 280 -525 300 -455
rect 215 -675 235 -605
rect 280 -675 300 -605
rect 200 -765 300 -745
rect 200 -830 300 -810
rect 200 -895 300 -875
rect 200 -960 300 -940
rect 225 -1040 295 -1020
rect 225 -1105 295 -1085
rect 225 -1170 295 -1150
rect 225 -1250 295 -1230
rect 225 -1315 295 -1295
rect 225 -1380 295 -1360
<< pdiffc >>
rect 225 380 295 400
rect 225 315 295 335
rect 225 250 295 270
rect 225 170 295 190
rect 225 105 295 125
rect 225 40 295 60
rect 215 -90 235 -20
rect 280 -90 300 -20
rect 215 -220 235 -150
rect 280 -220 300 -150
rect 215 -370 235 -300
rect 280 -370 300 -300
<< psubdiff >>
rect 90 -1305 140 -1290
rect 90 -1375 105 -1305
rect 125 -1375 140 -1305
rect 90 -1390 140 -1375
<< nsubdiff >>
rect 380 405 430 420
rect 380 335 395 405
rect 415 335 430 405
rect 380 320 430 335
<< psubdiffcont >>
rect 105 -1375 125 -1305
<< nsubdiffcont >>
rect 395 335 415 405
<< poly >>
rect 195 350 210 365
rect 310 355 365 365
rect 310 350 335 355
rect 325 335 335 350
rect 355 335 365 355
rect 325 325 365 335
rect 155 290 210 300
rect 155 270 165 290
rect 185 285 210 290
rect 310 285 405 300
rect 185 270 195 285
rect 155 260 195 270
rect 155 210 195 220
rect 155 190 165 210
rect 185 190 195 210
rect 155 180 195 190
rect 155 90 170 180
rect 195 140 210 155
rect 310 145 365 155
rect 310 140 335 145
rect 325 125 335 140
rect 355 125 365 145
rect 325 115 365 125
rect 155 75 210 90
rect 310 75 325 90
rect 105 -105 145 -95
rect 105 -125 115 -105
rect 135 -125 145 -105
rect 105 -135 145 -125
rect 105 -355 120 -135
rect 170 -230 185 75
rect 250 -5 265 10
rect 250 -135 265 -105
rect 145 -240 185 -230
rect 390 -180 405 285
rect 390 -195 410 -180
rect 145 -260 155 -240
rect 175 -260 185 -240
rect 145 -270 185 -260
rect 105 -365 145 -355
rect 105 -385 115 -365
rect 135 -385 145 -365
rect 105 -395 145 -385
rect 170 -445 185 -270
rect 250 -285 265 -235
rect 330 -240 370 -230
rect 330 -260 340 -240
rect 360 -260 370 -240
rect 330 -270 370 -260
rect 250 -440 265 -385
rect 145 -455 185 -445
rect 145 -475 155 -455
rect 175 -475 185 -455
rect 145 -485 185 -475
rect 170 -700 185 -485
rect 250 -590 265 -540
rect 335 -545 350 -270
rect 395 -280 410 -195
rect 390 -295 410 -280
rect 390 -330 405 -295
rect 390 -340 430 -330
rect 390 -360 400 -340
rect 420 -360 430 -340
rect 390 -370 430 -360
rect 325 -555 365 -545
rect 325 -575 335 -555
rect 355 -575 365 -555
rect 325 -585 365 -575
rect 130 -715 185 -700
rect 250 -705 265 -690
rect 130 -1060 145 -715
rect 250 -720 345 -705
rect 330 -780 345 -720
rect 170 -795 185 -780
rect 315 -795 345 -780
rect 330 -845 345 -795
rect 170 -860 185 -845
rect 315 -860 345 -845
rect 330 -910 345 -860
rect 170 -925 185 -910
rect 315 -925 450 -910
rect 115 -1075 145 -1060
rect 195 -1070 210 -1055
rect 310 -1070 365 -1055
rect 115 -1160 130 -1075
rect 155 -1105 195 -1095
rect 155 -1125 165 -1105
rect 185 -1120 195 -1105
rect 185 -1125 210 -1120
rect 155 -1135 210 -1125
rect 310 -1135 325 -1120
rect 115 -1175 170 -1160
rect 155 -1305 170 -1175
rect 350 -1160 365 -1070
rect 325 -1170 365 -1160
rect 325 -1190 335 -1170
rect 355 -1185 365 -1170
rect 355 -1190 410 -1185
rect 325 -1200 410 -1190
rect 325 -1250 365 -1240
rect 325 -1265 335 -1250
rect 195 -1280 210 -1265
rect 310 -1270 335 -1265
rect 355 -1270 365 -1250
rect 310 -1280 365 -1270
rect 155 -1315 195 -1305
rect 155 -1335 165 -1315
rect 185 -1330 195 -1315
rect 395 -1305 410 -1200
rect 370 -1315 410 -1305
rect 185 -1335 210 -1330
rect 155 -1345 210 -1335
rect 310 -1345 325 -1330
rect 370 -1335 380 -1315
rect 400 -1335 410 -1315
rect 370 -1345 410 -1335
rect 435 -1420 450 -925
rect 410 -1430 450 -1420
rect 410 -1450 420 -1430
rect 440 -1450 450 -1430
rect 410 -1460 450 -1450
<< polycont >>
rect 335 335 355 355
rect 165 270 185 290
rect 165 190 185 210
rect 335 125 355 145
rect 115 -125 135 -105
rect 155 -260 175 -240
rect 115 -385 135 -365
rect 340 -260 360 -240
rect 155 -475 175 -455
rect 400 -360 420 -340
rect 335 -575 355 -555
rect 165 -1125 185 -1105
rect 335 -1190 355 -1170
rect 335 -1270 355 -1250
rect 165 -1335 185 -1315
rect 380 -1335 400 -1315
rect 420 -1450 440 -1430
<< locali >>
rect 215 400 305 410
rect 215 390 225 400
rect 165 380 225 390
rect 295 380 305 400
rect 165 370 305 380
rect 385 405 425 415
rect 165 300 185 370
rect 325 355 365 365
rect 215 335 305 345
rect 215 315 225 335
rect 295 315 305 335
rect 325 335 335 355
rect 355 335 365 355
rect 325 325 365 335
rect 385 335 395 405
rect 415 335 425 405
rect 385 325 425 335
rect 215 305 305 315
rect 155 290 195 300
rect 155 280 165 290
rect 115 270 165 280
rect 185 270 195 290
rect 115 260 195 270
rect 215 270 305 280
rect 115 -95 135 260
rect 215 250 225 270
rect 295 260 305 270
rect 330 260 350 325
rect 295 250 390 260
rect 215 240 390 250
rect 155 210 195 220
rect 155 190 165 210
rect 185 200 195 210
rect 185 190 305 200
rect 155 180 225 190
rect 215 170 225 180
rect 295 170 305 190
rect 370 195 390 240
rect 370 175 405 195
rect 215 160 305 170
rect 325 145 365 155
rect 215 125 305 135
rect 215 115 225 125
rect 175 105 225 115
rect 295 105 305 125
rect 325 125 335 145
rect 355 125 365 145
rect 325 115 365 125
rect 175 95 305 105
rect 175 -10 195 95
rect 215 60 305 70
rect 215 40 225 60
rect 295 50 305 60
rect 330 50 350 115
rect 385 95 405 175
rect 295 40 350 50
rect 215 30 350 40
rect 175 -20 245 -10
rect 175 -30 215 -20
rect 205 -90 215 -30
rect 235 -90 245 -20
rect 105 -105 145 -95
rect 205 -100 245 -90
rect 270 -20 310 -10
rect 270 -90 280 -20
rect 300 -90 310 -20
rect 270 -100 310 -90
rect 105 -125 115 -105
rect 135 -125 145 -105
rect 105 -135 145 -125
rect 205 -150 245 -140
rect 205 -155 215 -150
rect 85 -175 215 -155
rect 205 -220 215 -175
rect 235 -220 245 -150
rect 205 -230 245 -220
rect 270 -150 310 -140
rect 270 -220 280 -150
rect 300 -220 310 -150
rect 270 -230 310 -220
rect 330 -230 350 30
rect 370 75 405 95
rect 370 -150 390 75
rect 370 -155 450 -150
rect 370 -170 470 -155
rect 370 -190 390 -170
rect 430 -175 470 -170
rect 370 -210 410 -190
rect 145 -240 185 -230
rect 145 -260 155 -240
rect 175 -250 185 -240
rect 270 -250 290 -230
rect 330 -240 370 -230
rect 330 -250 340 -240
rect 175 -260 290 -250
rect 145 -270 290 -260
rect 310 -260 340 -250
rect 360 -260 370 -240
rect 310 -270 370 -260
rect 310 -290 330 -270
rect 390 -290 410 -210
rect 205 -300 245 -290
rect 205 -315 215 -300
rect 85 -335 215 -315
rect 105 -365 145 -355
rect 105 -385 115 -365
rect 135 -385 145 -365
rect 205 -370 215 -335
rect 235 -370 245 -300
rect 205 -380 245 -370
rect 270 -300 330 -290
rect 270 -370 280 -300
rect 300 -310 330 -300
rect 350 -310 410 -290
rect 300 -370 310 -310
rect 270 -380 310 -370
rect 105 -395 145 -385
rect 105 -500 125 -395
rect 350 -445 370 -310
rect 430 -330 470 -315
rect 390 -335 470 -330
rect 390 -340 450 -335
rect 390 -360 400 -340
rect 420 -350 450 -340
rect 420 -360 430 -350
rect 390 -370 430 -360
rect 145 -455 245 -445
rect 145 -475 155 -455
rect 175 -465 215 -455
rect 175 -475 185 -465
rect 145 -485 185 -475
rect 105 -520 135 -500
rect 115 -665 135 -520
rect 205 -525 215 -465
rect 235 -525 245 -455
rect 205 -535 245 -525
rect 270 -455 390 -445
rect 270 -525 280 -455
rect 300 -465 390 -455
rect 300 -525 310 -465
rect 370 -505 390 -465
rect 370 -525 405 -505
rect 270 -535 310 -525
rect 325 -555 365 -545
rect 325 -575 335 -555
rect 355 -575 365 -555
rect 325 -585 365 -575
rect 205 -605 245 -595
rect 205 -665 215 -605
rect 115 -675 215 -665
rect 235 -675 245 -605
rect 115 -685 245 -675
rect 270 -605 310 -595
rect 330 -605 350 -585
rect 270 -675 280 -605
rect 300 -625 350 -605
rect 300 -675 310 -625
rect 270 -685 310 -675
rect 330 -670 350 -625
rect 385 -630 405 -525
rect 385 -650 435 -630
rect 115 -1030 135 -685
rect 330 -690 395 -670
rect 190 -745 310 -735
rect 190 -765 200 -745
rect 300 -765 310 -745
rect 190 -775 310 -765
rect 190 -810 310 -800
rect 190 -830 200 -810
rect 300 -820 310 -810
rect 300 -830 350 -820
rect 190 -840 350 -830
rect 190 -875 310 -865
rect 190 -895 200 -875
rect 300 -895 310 -875
rect 190 -905 310 -895
rect 330 -930 350 -840
rect 190 -940 350 -930
rect 190 -960 200 -940
rect 300 -950 350 -940
rect 300 -960 310 -950
rect 190 -970 310 -960
rect 215 -1020 305 -1010
rect 215 -1030 225 -1020
rect 115 -1040 225 -1030
rect 295 -1040 305 -1020
rect 115 -1050 305 -1040
rect 165 -1095 185 -1050
rect 330 -1075 350 -950
rect 215 -1085 350 -1075
rect 155 -1105 195 -1095
rect 155 -1125 165 -1105
rect 185 -1125 195 -1105
rect 215 -1105 225 -1085
rect 295 -1095 350 -1085
rect 295 -1105 305 -1095
rect 215 -1115 305 -1105
rect 155 -1135 195 -1125
rect 375 -1125 395 -690
rect 415 -1090 435 -650
rect 415 -1110 445 -1090
rect 215 -1150 305 -1140
rect 375 -1145 405 -1125
rect 215 -1170 225 -1150
rect 295 -1160 305 -1150
rect 295 -1170 365 -1160
rect 215 -1180 335 -1170
rect 325 -1190 335 -1180
rect 355 -1190 365 -1170
rect 325 -1200 365 -1190
rect 385 -1220 405 -1145
rect 215 -1230 305 -1220
rect 215 -1240 225 -1230
rect 165 -1250 225 -1240
rect 295 -1250 305 -1230
rect 375 -1240 405 -1220
rect 165 -1260 305 -1250
rect 325 -1250 395 -1240
rect 95 -1305 135 -1295
rect 165 -1305 185 -1260
rect 325 -1270 335 -1250
rect 355 -1260 395 -1250
rect 355 -1270 365 -1260
rect 325 -1280 365 -1270
rect 215 -1295 305 -1285
rect 95 -1375 105 -1305
rect 125 -1375 135 -1305
rect 155 -1315 195 -1305
rect 155 -1335 165 -1315
rect 185 -1335 195 -1315
rect 215 -1315 225 -1295
rect 295 -1315 305 -1295
rect 215 -1325 305 -1315
rect 155 -1345 195 -1335
rect 330 -1350 350 -1280
rect 425 -1305 445 -1110
rect 370 -1315 445 -1305
rect 370 -1335 380 -1315
rect 400 -1325 445 -1315
rect 400 -1335 410 -1325
rect 370 -1345 410 -1335
rect 95 -1385 135 -1375
rect 215 -1360 350 -1350
rect 215 -1380 225 -1360
rect 295 -1370 350 -1360
rect 295 -1380 305 -1370
rect 215 -1390 305 -1380
rect 410 -1430 450 -1420
rect 410 -1450 420 -1430
rect 440 -1450 450 -1430
rect 410 -1460 450 -1450
<< viali >>
rect 225 315 295 335
rect 395 335 415 405
rect 280 -90 300 -20
rect 200 -765 300 -745
rect 200 -895 300 -875
rect 105 -1375 125 -1305
rect 225 -1315 295 -1295
rect 420 -1450 440 -1430
<< metal1 >>
rect 85 405 470 420
rect 85 335 395 405
rect 415 335 470 405
rect 85 315 225 335
rect 295 315 470 335
rect 85 -20 470 315
rect 85 -90 280 -20
rect 300 -90 470 -20
rect 85 -105 470 -90
rect 85 -745 470 -730
rect 85 -765 200 -745
rect 300 -765 470 -745
rect 85 -875 470 -765
rect 85 -895 200 -875
rect 300 -895 470 -875
rect 85 -1295 470 -895
rect 85 -1305 225 -1295
rect 85 -1375 105 -1305
rect 125 -1315 225 -1305
rect 295 -1315 470 -1295
rect 125 -1375 470 -1315
rect 85 -1390 470 -1375
rect 85 -1430 470 -1420
rect 85 -1450 420 -1430
rect 440 -1450 470 -1430
rect 85 -1460 470 -1450
<< labels >>
rlabel locali 85 -165 85 -165 7 D
rlabel locali 85 -325 85 -325 7 D_BAR
rlabel locali 470 -165 470 -165 3 Q
rlabel locali 470 -325 470 -325 3 Q_BAR
rlabel metal1 85 155 85 155 7 VP
rlabel metal1 85 -1270 85 -1270 7 VN
rlabel metal1 85 -1440 85 -1440 7 CLK
<< end >>
