magic
tech sky130A
timestamp 1695761726
<< nwell >>
rect -85 -345 230 545
<< nmos >>
rect 20 -460 120 -445
rect 20 -605 120 -590
rect 40 -1060 55 -690
rect 20 -1190 120 -1175
rect 20 -1255 120 -1240
rect 20 -1400 120 -1385
rect 20 -1465 120 -1450
<< pmos >>
rect 20 460 120 475
rect 20 395 120 410
rect 20 250 120 265
rect 20 185 120 200
rect 20 15 120 30
rect 20 -130 120 -115
rect 20 -275 120 -260
<< ndiff >>
rect 20 -410 120 -395
rect 20 -430 35 -410
rect 105 -430 120 -410
rect 20 -445 120 -430
rect 20 -475 120 -460
rect 20 -495 35 -475
rect 105 -495 120 -475
rect 20 -510 120 -495
rect 20 -555 120 -540
rect 20 -575 35 -555
rect 105 -575 120 -555
rect 20 -590 120 -575
rect 20 -620 120 -605
rect 20 -640 35 -620
rect 105 -640 120 -620
rect 20 -655 120 -640
rect -10 -705 40 -690
rect -10 -1045 5 -705
rect 25 -1045 40 -705
rect -10 -1060 40 -1045
rect 55 -705 105 -690
rect 55 -1045 70 -705
rect 90 -1045 105 -705
rect 55 -1060 105 -1045
rect 20 -1140 120 -1125
rect 20 -1160 35 -1140
rect 105 -1160 120 -1140
rect 20 -1175 120 -1160
rect 20 -1205 120 -1190
rect 20 -1225 35 -1205
rect 105 -1225 120 -1205
rect 20 -1240 120 -1225
rect 20 -1270 120 -1255
rect 20 -1290 35 -1270
rect 105 -1290 120 -1270
rect 20 -1305 120 -1290
rect 20 -1350 120 -1335
rect 20 -1370 35 -1350
rect 105 -1370 120 -1350
rect 20 -1385 120 -1370
rect 20 -1415 120 -1400
rect 20 -1435 35 -1415
rect 105 -1435 120 -1415
rect 20 -1450 120 -1435
rect 20 -1480 120 -1465
rect 20 -1500 35 -1480
rect 105 -1500 120 -1480
rect 20 -1515 120 -1500
<< pdiff >>
rect 20 510 120 525
rect 20 490 35 510
rect 105 490 120 510
rect 20 475 120 490
rect 20 445 120 460
rect 20 425 35 445
rect 105 425 120 445
rect 20 410 120 425
rect 20 380 120 395
rect 20 360 35 380
rect 105 360 120 380
rect 20 345 120 360
rect 20 300 120 315
rect 20 280 35 300
rect 105 280 120 300
rect 20 265 120 280
rect 20 235 120 250
rect 20 215 35 235
rect 105 215 120 235
rect 20 200 120 215
rect 20 170 120 185
rect 20 150 35 170
rect 105 150 120 170
rect 20 135 120 150
rect 20 65 120 80
rect 20 45 35 65
rect 105 45 120 65
rect 20 30 120 45
rect 20 0 120 15
rect 20 -20 35 0
rect 105 -20 120 0
rect 20 -35 120 -20
rect 20 -80 120 -65
rect 20 -100 35 -80
rect 105 -100 120 -80
rect 20 -115 120 -100
rect 20 -145 120 -130
rect 20 -165 35 -145
rect 105 -165 120 -145
rect 20 -180 120 -165
rect 20 -225 120 -210
rect 20 -245 35 -225
rect 105 -245 120 -225
rect 20 -260 120 -245
rect 20 -290 120 -275
rect 20 -310 35 -290
rect 105 -310 120 -290
rect 20 -325 120 -310
<< ndiffc >>
rect 35 -430 105 -410
rect 35 -495 105 -475
rect 35 -575 105 -555
rect 35 -640 105 -620
rect 5 -1045 25 -705
rect 70 -1045 90 -705
rect 35 -1160 105 -1140
rect 35 -1225 105 -1205
rect 35 -1290 105 -1270
rect 35 -1370 105 -1350
rect 35 -1435 105 -1415
rect 35 -1500 105 -1480
<< pdiffc >>
rect 35 490 105 510
rect 35 425 105 445
rect 35 360 105 380
rect 35 280 105 300
rect 35 215 105 235
rect 35 150 105 170
rect 35 45 105 65
rect 35 -20 105 0
rect 35 -100 105 -80
rect 35 -165 105 -145
rect 35 -245 105 -225
rect 35 -310 105 -290
<< psubdiff >>
rect -60 -1330 -10 -1315
rect -60 -1400 -45 -1330
rect -25 -1400 -10 -1330
rect -60 -1415 -10 -1400
<< nsubdiff >>
rect 150 390 200 405
rect 150 320 165 390
rect 185 320 200 390
rect 150 305 200 320
<< psubdiffcont >>
rect -45 -1400 -25 -1330
<< nsubdiffcont >>
rect 165 320 185 390
<< poly >>
rect -75 460 20 475
rect 120 460 135 475
rect -75 370 -60 460
rect -35 425 5 435
rect -35 405 -25 425
rect -5 410 5 425
rect -5 405 20 410
rect -35 395 20 405
rect 120 395 135 410
rect -75 360 -35 370
rect -75 340 -65 360
rect -45 340 -35 360
rect -75 330 -35 340
rect -75 -340 -60 330
rect -10 305 5 395
rect -35 290 5 305
rect -35 -50 -20 290
rect 5 250 20 265
rect 120 250 215 265
rect 135 215 175 225
rect 135 200 145 215
rect 5 185 20 200
rect 120 195 145 200
rect 165 195 175 215
rect 120 185 175 195
rect 135 95 150 185
rect 200 160 215 250
rect 175 150 215 160
rect 175 130 185 150
rect 205 130 215 150
rect 175 120 215 130
rect 135 85 175 95
rect 135 65 145 85
rect 165 65 175 85
rect 135 55 175 65
rect 200 30 215 120
rect 5 15 20 30
rect 120 15 145 30
rect -35 -60 5 -50
rect -35 -80 -25 -60
rect -5 -80 5 -60
rect -35 -90 5 -80
rect -35 -300 -20 -90
rect 130 -115 145 15
rect 5 -130 20 -115
rect 120 -130 145 -115
rect 130 -260 145 -130
rect 5 -275 20 -260
rect 120 -275 145 -260
rect -35 -315 5 -300
rect -75 -350 -35 -340
rect -75 -370 -65 -350
rect -45 -370 -35 -350
rect -75 -380 -35 -370
rect -75 -1110 -60 -380
rect -10 -405 5 -315
rect 130 -340 145 -275
rect 50 -350 145 -340
rect 50 -370 60 -350
rect 80 -355 145 -350
rect 80 -370 90 -355
rect 50 -380 90 -370
rect -35 -420 5 -405
rect -35 -525 -20 -420
rect 130 -445 145 -355
rect 5 -460 20 -445
rect 120 -460 145 -445
rect -35 -535 5 -525
rect -35 -555 -25 -535
rect -5 -555 5 -535
rect -35 -565 5 -555
rect -35 -1070 -20 -565
rect 130 -590 145 -460
rect 5 -605 20 -590
rect 120 -605 145 -590
rect 130 -665 145 -605
rect 40 -680 145 -665
rect 170 15 215 30
rect 40 -690 55 -680
rect 170 -705 185 15
rect 120 -715 185 -705
rect 120 -735 130 -715
rect 150 -720 185 -715
rect 150 -735 160 -720
rect 120 -745 160 -735
rect -35 -1085 5 -1070
rect 40 -1075 55 -1060
rect -75 -1120 -35 -1110
rect -75 -1140 -65 -1120
rect -45 -1140 -35 -1120
rect -75 -1150 -35 -1140
rect -75 -1240 -60 -1150
rect -10 -1175 5 -1085
rect 120 -1100 135 -745
rect 160 -780 200 -770
rect 160 -800 170 -780
rect 190 -800 200 -780
rect 160 -810 200 -800
rect 160 -1060 175 -810
rect 160 -1075 215 -1060
rect 120 -1115 175 -1100
rect -35 -1185 20 -1175
rect -35 -1205 -25 -1185
rect -5 -1190 20 -1185
rect 120 -1190 135 -1175
rect -5 -1205 5 -1190
rect -35 -1215 5 -1205
rect -75 -1255 20 -1240
rect 120 -1255 135 -1240
rect 160 -1280 175 -1115
rect 135 -1295 175 -1280
rect 135 -1385 150 -1295
rect 200 -1320 215 -1075
rect 175 -1330 215 -1320
rect 175 -1350 185 -1330
rect 205 -1350 215 -1330
rect 175 -1360 215 -1350
rect 5 -1400 20 -1385
rect 120 -1395 175 -1385
rect 120 -1400 145 -1395
rect 135 -1415 145 -1400
rect 165 -1415 175 -1395
rect 135 -1425 175 -1415
rect 200 -1450 215 -1360
rect 5 -1465 20 -1450
rect 120 -1465 215 -1450
<< polycont >>
rect -25 405 -5 425
rect -65 340 -45 360
rect 145 195 165 215
rect 185 130 205 150
rect 145 65 165 85
rect -25 -80 -5 -60
rect -65 -370 -45 -350
rect 60 -370 80 -350
rect -25 -555 -5 -535
rect 130 -735 150 -715
rect -65 -1140 -45 -1120
rect 170 -800 190 -780
rect -25 -1205 -5 -1185
rect 185 -1350 205 -1330
rect 145 -1415 165 -1395
<< locali >>
rect -15 510 115 520
rect -15 500 35 510
rect -15 435 5 500
rect 25 490 35 500
rect 105 490 115 510
rect 25 480 115 490
rect -35 425 5 435
rect -35 405 -25 425
rect -5 405 5 425
rect 25 445 115 455
rect 25 425 35 445
rect 105 425 115 445
rect 25 415 115 425
rect -35 395 5 405
rect 155 390 195 400
rect 25 380 115 390
rect 25 370 35 380
rect -75 360 35 370
rect 105 360 115 380
rect -75 340 -65 360
rect -45 350 115 360
rect -45 340 -35 350
rect -75 330 -35 340
rect 155 320 165 390
rect 185 320 195 390
rect 155 310 195 320
rect 25 300 115 310
rect 25 280 35 300
rect 105 290 115 300
rect 105 280 155 290
rect 25 270 155 280
rect 25 235 115 245
rect 25 225 35 235
rect -15 215 35 225
rect 105 215 115 235
rect -15 205 115 215
rect 135 225 155 270
rect 135 215 175 225
rect -15 75 5 205
rect 135 195 145 215
rect 165 195 175 215
rect 135 185 175 195
rect 25 170 115 180
rect 25 150 35 170
rect 105 160 115 170
rect 105 150 215 160
rect 25 140 185 150
rect 175 130 185 140
rect 205 130 215 150
rect 175 120 215 130
rect 135 85 175 95
rect -15 65 115 75
rect -15 55 35 65
rect 25 45 35 55
rect 105 45 115 65
rect 135 65 145 85
rect 165 65 175 85
rect 135 55 175 65
rect 25 35 115 45
rect 25 0 115 10
rect 25 -20 35 0
rect 105 -20 115 0
rect 25 -30 115 -20
rect -35 -60 5 -50
rect -35 -80 -25 -60
rect -5 -70 5 -60
rect -5 -80 115 -70
rect -35 -90 35 -80
rect 25 -100 35 -90
rect 105 -100 115 -80
rect 25 -110 115 -100
rect 25 -145 115 -135
rect 25 -155 35 -145
rect -85 -165 35 -155
rect 105 -165 115 -145
rect -85 -175 115 -165
rect 140 -215 160 55
rect 195 -155 215 120
rect 195 -175 230 -155
rect -85 -225 115 -215
rect -85 -235 35 -225
rect 25 -245 35 -235
rect 105 -245 115 -225
rect 25 -255 115 -245
rect 140 -235 230 -215
rect 25 -290 115 -280
rect 25 -300 35 -290
rect -55 -310 35 -300
rect 105 -310 115 -290
rect -55 -320 115 -310
rect -55 -340 -35 -320
rect -75 -350 -35 -340
rect -75 -370 -65 -350
rect -45 -370 -35 -350
rect -75 -380 -35 -370
rect 50 -350 90 -340
rect 50 -370 60 -350
rect 80 -370 90 -350
rect 50 -380 90 -370
rect -55 -400 -35 -380
rect -55 -410 115 -400
rect -55 -420 35 -410
rect 25 -430 35 -420
rect 105 -430 115 -410
rect 25 -440 115 -430
rect 140 -465 160 -235
rect 25 -475 160 -465
rect 25 -495 35 -475
rect 105 -485 160 -475
rect 105 -495 115 -485
rect 25 -505 115 -495
rect -35 -535 5 -525
rect -35 -555 -25 -535
rect -5 -545 5 -535
rect -5 -555 115 -545
rect -35 -565 35 -555
rect 25 -575 35 -565
rect 105 -575 115 -555
rect 25 -585 115 -575
rect 140 -590 160 -485
rect 140 -610 200 -590
rect 25 -620 115 -610
rect 25 -640 35 -620
rect 105 -630 115 -620
rect 105 -640 140 -630
rect 25 -650 140 -640
rect -5 -705 35 -695
rect -5 -1045 5 -705
rect 25 -1045 35 -705
rect -5 -1055 35 -1045
rect 60 -705 100 -695
rect 60 -1045 70 -705
rect 90 -1045 100 -705
rect 120 -705 140 -650
rect 120 -715 160 -705
rect 120 -735 130 -715
rect 150 -735 160 -715
rect 120 -745 160 -735
rect 180 -770 200 -610
rect 160 -780 200 -770
rect 160 -800 170 -780
rect 190 -800 200 -780
rect 160 -810 200 -800
rect 60 -1055 100 -1045
rect 80 -1090 100 -1055
rect 80 -1110 155 -1090
rect -75 -1120 -35 -1110
rect -75 -1140 -65 -1120
rect -45 -1130 -35 -1120
rect -45 -1140 115 -1130
rect -75 -1150 35 -1140
rect 25 -1160 35 -1150
rect 105 -1160 115 -1140
rect 25 -1170 115 -1160
rect -35 -1185 5 -1175
rect -35 -1205 -25 -1185
rect -5 -1205 5 -1185
rect 135 -1195 155 -1110
rect -35 -1215 5 -1205
rect -15 -1280 5 -1215
rect 25 -1205 155 -1195
rect 25 -1225 35 -1205
rect 105 -1215 155 -1205
rect 105 -1225 115 -1215
rect 25 -1235 115 -1225
rect 25 -1270 115 -1260
rect 25 -1280 35 -1270
rect -15 -1290 35 -1280
rect 105 -1290 115 -1270
rect -15 -1300 115 -1290
rect -55 -1330 -15 -1320
rect -55 -1400 -45 -1330
rect -25 -1400 -15 -1330
rect 175 -1330 215 -1320
rect 175 -1340 185 -1330
rect 25 -1350 185 -1340
rect 205 -1350 215 -1330
rect 25 -1370 35 -1350
rect 105 -1360 215 -1350
rect 105 -1370 115 -1360
rect 25 -1380 115 -1370
rect -55 -1410 -15 -1400
rect 135 -1395 175 -1385
rect 25 -1415 115 -1405
rect 25 -1435 35 -1415
rect 105 -1435 115 -1415
rect 25 -1445 115 -1435
rect 135 -1415 145 -1395
rect 165 -1415 175 -1395
rect 135 -1425 175 -1415
rect 135 -1470 155 -1425
rect 25 -1480 155 -1470
rect 25 -1500 35 -1480
rect 105 -1490 155 -1480
rect 105 -1500 115 -1490
rect 25 -1510 115 -1500
<< viali >>
rect 35 425 105 445
rect 165 320 185 390
rect 35 -20 105 0
rect 5 -1045 25 -705
rect -45 -1400 -25 -1330
rect 35 -1435 105 -1415
<< metal1 >>
rect -85 445 230 460
rect -85 425 35 445
rect 105 425 230 445
rect -85 390 230 425
rect -85 320 165 390
rect 185 320 230 390
rect -85 0 230 320
rect -85 -20 35 0
rect 105 -20 230 0
rect -85 -35 230 -20
rect -85 -380 230 -340
rect -85 -705 230 -690
rect -85 -1045 5 -705
rect 25 -1045 230 -705
rect -85 -1330 230 -1045
rect -85 -1400 -45 -1330
rect -25 -1400 230 -1330
rect -85 -1415 230 -1400
rect -85 -1435 35 -1415
rect 105 -1435 230 -1415
rect -85 -1450 230 -1435
<< end >>
