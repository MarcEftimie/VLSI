magic
tech sky130A
timestamp 1697389219
<< nwell >>
rect 550 -1180 4140 205
<< nmos >>
rect 845 -2455 895 -1255
rect 1075 -2455 1125 -1255
rect 1175 -2455 1225 -1255
rect 1275 -2455 1325 -1255
rect 1375 -2455 1425 -1255
rect 1475 -2455 1525 -1255
rect 1575 -2455 1625 -1255
rect 1675 -2455 1725 -1255
rect 1775 -2455 1825 -1255
rect 1875 -2455 1925 -1255
rect 1975 -2455 2025 -1255
rect 2075 -2455 2125 -1255
rect 2175 -2455 2225 -1255
rect 2275 -2455 2325 -1255
rect 2375 -2455 2425 -1255
rect 2670 -2455 2720 -1255
rect 2770 -2455 2820 -1255
rect 2870 -2455 2920 -1255
rect 2970 -2455 3020 -1255
rect 3070 -2455 3120 -1255
rect 3170 -2455 3220 -1255
rect 3270 -2455 3320 -1255
rect 3370 -2455 3420 -1255
rect 3470 -2455 3520 -1255
rect 3570 -2455 3620 -1255
rect 3670 -2455 3720 -1255
rect 3770 -2455 3820 -1255
rect 3870 -2455 3920 -1255
rect 3970 -2455 4020 -1255
<< pmos >>
rect 605 0 905 50
rect 605 -100 905 -50
rect 605 -200 905 -150
rect 605 -300 905 -250
rect 605 -400 905 -350
rect 605 -500 905 -450
rect 605 -600 905 -550
rect 605 -700 905 -650
rect 605 -800 905 -750
rect 605 -900 905 -850
rect 1075 -1055 1125 145
rect 1175 -1055 1225 145
rect 1275 -1055 1325 145
rect 1375 -1055 1425 145
rect 1475 -1055 1525 145
rect 1575 -1055 1625 145
rect 1675 -1055 1725 145
rect 1775 -1055 1825 145
rect 1875 -1055 1925 145
rect 1975 -1055 2025 145
rect 2075 -1055 2125 145
rect 2175 -1055 2225 145
rect 2275 -1055 2325 145
rect 2375 -1055 2425 145
rect 2670 -1120 2720 80
rect 2770 -1120 2820 80
rect 2870 -1120 2920 80
rect 2970 -1120 3020 80
rect 3070 -1120 3120 80
rect 3170 -1120 3220 80
rect 3270 -1120 3320 80
rect 3370 -1120 3420 80
rect 3470 -1120 3520 80
rect 3570 -1120 3620 80
rect 3670 -1120 3720 80
rect 3770 -1120 3820 80
rect 3870 -1120 3920 80
rect 3970 -1120 4020 80
<< ndiff >>
rect 795 -1270 845 -1255
rect 795 -2435 810 -1270
rect 830 -2435 845 -1270
rect 795 -2455 845 -2435
rect 895 -1270 945 -1255
rect 895 -2435 910 -1270
rect 930 -2435 945 -1270
rect 895 -2455 945 -2435
rect 1025 -1270 1075 -1255
rect 1025 -2440 1040 -1270
rect 1060 -2440 1075 -1270
rect 1025 -2455 1075 -2440
rect 1125 -1270 1175 -1255
rect 1125 -2440 1140 -1270
rect 1160 -2440 1175 -1270
rect 1125 -2455 1175 -2440
rect 1225 -1270 1275 -1255
rect 1225 -2440 1240 -1270
rect 1260 -2440 1275 -1270
rect 1225 -2455 1275 -2440
rect 1325 -1270 1375 -1255
rect 1325 -2440 1340 -1270
rect 1360 -2440 1375 -1270
rect 1325 -2455 1375 -2440
rect 1425 -1270 1475 -1255
rect 1425 -2440 1440 -1270
rect 1460 -2440 1475 -1270
rect 1425 -2455 1475 -2440
rect 1525 -1270 1575 -1255
rect 1525 -2440 1540 -1270
rect 1560 -2440 1575 -1270
rect 1525 -2455 1575 -2440
rect 1625 -1270 1675 -1255
rect 1625 -2440 1640 -1270
rect 1660 -2440 1675 -1270
rect 1625 -2455 1675 -2440
rect 1725 -1270 1775 -1255
rect 1725 -2440 1740 -1270
rect 1760 -2440 1775 -1270
rect 1725 -2455 1775 -2440
rect 1825 -1270 1875 -1255
rect 1825 -2440 1840 -1270
rect 1860 -2440 1875 -1270
rect 1825 -2455 1875 -2440
rect 1925 -1270 1975 -1255
rect 1925 -2440 1940 -1270
rect 1960 -2440 1975 -1270
rect 1925 -2455 1975 -2440
rect 2025 -1270 2075 -1255
rect 2025 -2440 2040 -1270
rect 2060 -2440 2075 -1270
rect 2025 -2455 2075 -2440
rect 2125 -1270 2175 -1255
rect 2125 -2440 2140 -1270
rect 2160 -2440 2175 -1270
rect 2125 -2455 2175 -2440
rect 2225 -1270 2275 -1255
rect 2225 -2440 2240 -1270
rect 2260 -2440 2275 -1270
rect 2225 -2455 2275 -2440
rect 2325 -1270 2375 -1255
rect 2325 -2440 2340 -1270
rect 2360 -2440 2375 -1270
rect 2325 -2455 2375 -2440
rect 2425 -1270 2470 -1255
rect 2425 -2440 2440 -1270
rect 2460 -2440 2470 -1270
rect 2425 -2455 2470 -2440
rect 2625 -1270 2670 -1255
rect 2625 -2440 2635 -1270
rect 2655 -2440 2670 -1270
rect 2625 -2455 2670 -2440
rect 2720 -1270 2770 -1255
rect 2720 -2440 2735 -1270
rect 2755 -2440 2770 -1270
rect 2720 -2455 2770 -2440
rect 2820 -1270 2870 -1255
rect 2820 -2440 2835 -1270
rect 2855 -2440 2870 -1270
rect 2820 -2455 2870 -2440
rect 2920 -1270 2970 -1255
rect 2920 -2440 2935 -1270
rect 2955 -2440 2970 -1270
rect 2920 -2455 2970 -2440
rect 3020 -1270 3070 -1255
rect 3020 -2440 3035 -1270
rect 3055 -2440 3070 -1270
rect 3020 -2455 3070 -2440
rect 3120 -1270 3170 -1255
rect 3120 -2440 3135 -1270
rect 3155 -2440 3170 -1270
rect 3120 -2455 3170 -2440
rect 3220 -1270 3270 -1255
rect 3220 -2440 3235 -1270
rect 3255 -2440 3270 -1270
rect 3220 -2455 3270 -2440
rect 3320 -1270 3370 -1255
rect 3320 -2440 3335 -1270
rect 3355 -2440 3370 -1270
rect 3320 -2455 3370 -2440
rect 3420 -1270 3470 -1255
rect 3420 -2440 3435 -1270
rect 3455 -2440 3470 -1270
rect 3420 -2455 3470 -2440
rect 3520 -1270 3570 -1255
rect 3520 -2440 3535 -1270
rect 3555 -2440 3570 -1270
rect 3520 -2455 3570 -2440
rect 3620 -1270 3670 -1255
rect 3620 -2440 3635 -1270
rect 3655 -2440 3670 -1270
rect 3620 -2455 3670 -2440
rect 3720 -1270 3770 -1255
rect 3720 -2440 3735 -1270
rect 3755 -2440 3770 -1270
rect 3720 -2455 3770 -2440
rect 3820 -1270 3870 -1255
rect 3820 -2440 3835 -1270
rect 3855 -2440 3870 -1270
rect 3820 -2455 3870 -2440
rect 3920 -1270 3970 -1255
rect 3920 -2440 3935 -1270
rect 3955 -2440 3970 -1270
rect 3920 -2455 3970 -2440
rect 4020 -1270 4070 -1255
rect 4020 -2440 4035 -1270
rect 4055 -2440 4070 -1270
rect 4020 -2455 4070 -2440
<< pdiff >>
rect 605 85 905 95
rect 605 65 620 85
rect 890 65 905 85
rect 605 50 905 65
rect 1025 130 1075 145
rect 605 -15 905 0
rect 605 -35 620 -15
rect 890 -35 905 -15
rect 605 -50 905 -35
rect 605 -115 905 -100
rect 605 -135 620 -115
rect 890 -135 905 -115
rect 605 -150 905 -135
rect 605 -215 905 -200
rect 605 -235 620 -215
rect 890 -235 905 -215
rect 605 -250 905 -235
rect 605 -315 905 -300
rect 605 -335 620 -315
rect 890 -335 905 -315
rect 605 -350 905 -335
rect 605 -415 905 -400
rect 605 -435 620 -415
rect 890 -435 905 -415
rect 605 -450 905 -435
rect 605 -515 905 -500
rect 605 -535 620 -515
rect 890 -535 905 -515
rect 605 -550 905 -535
rect 605 -615 905 -600
rect 605 -635 620 -615
rect 890 -635 905 -615
rect 605 -650 905 -635
rect 605 -715 905 -700
rect 605 -735 620 -715
rect 890 -735 905 -715
rect 605 -750 905 -735
rect 605 -815 905 -800
rect 605 -835 620 -815
rect 890 -835 905 -815
rect 605 -850 905 -835
rect 605 -915 905 -900
rect 605 -935 620 -915
rect 890 -935 905 -915
rect 605 -950 905 -935
rect 1025 -1040 1040 130
rect 1060 -1040 1075 130
rect 1025 -1055 1075 -1040
rect 1125 130 1175 145
rect 1125 -1040 1140 130
rect 1160 -1040 1175 130
rect 1125 -1055 1175 -1040
rect 1225 130 1275 145
rect 1225 -1040 1240 130
rect 1260 -1040 1275 130
rect 1225 -1055 1275 -1040
rect 1325 130 1375 145
rect 1325 -1040 1340 130
rect 1360 -1040 1375 130
rect 1325 -1055 1375 -1040
rect 1425 130 1475 145
rect 1425 -1040 1440 130
rect 1460 -1040 1475 130
rect 1425 -1055 1475 -1040
rect 1525 130 1575 145
rect 1525 -1040 1540 130
rect 1560 -1040 1575 130
rect 1525 -1055 1575 -1040
rect 1625 130 1675 145
rect 1625 -1040 1640 130
rect 1660 -1040 1675 130
rect 1625 -1055 1675 -1040
rect 1725 130 1775 145
rect 1725 -1040 1740 130
rect 1760 -1040 1775 130
rect 1725 -1055 1775 -1040
rect 1825 130 1875 145
rect 1825 -1040 1840 130
rect 1860 -1040 1875 130
rect 1825 -1055 1875 -1040
rect 1925 130 1975 145
rect 1925 -1040 1940 130
rect 1960 -1040 1975 130
rect 1925 -1055 1975 -1040
rect 2025 130 2075 145
rect 2025 -1040 2040 130
rect 2060 -1040 2075 130
rect 2025 -1055 2075 -1040
rect 2125 130 2175 145
rect 2125 -1040 2140 130
rect 2160 -1040 2175 130
rect 2125 -1055 2175 -1040
rect 2225 130 2275 145
rect 2225 -1040 2240 130
rect 2260 -1040 2275 130
rect 2225 -1055 2275 -1040
rect 2325 130 2375 145
rect 2325 -1040 2340 130
rect 2360 -1040 2375 130
rect 2325 -1055 2375 -1040
rect 2425 130 2470 145
rect 2425 -1040 2440 130
rect 2460 -1040 2470 130
rect 2425 -1055 2470 -1040
rect 2625 65 2670 80
rect 2625 -1105 2635 65
rect 2655 -1105 2670 65
rect 2625 -1120 2670 -1105
rect 2720 65 2770 80
rect 2720 -1105 2735 65
rect 2755 -1105 2770 65
rect 2720 -1120 2770 -1105
rect 2820 65 2870 80
rect 2820 -1105 2835 65
rect 2855 -1105 2870 65
rect 2820 -1120 2870 -1105
rect 2920 65 2970 80
rect 2920 -1105 2935 65
rect 2955 -1105 2970 65
rect 2920 -1120 2970 -1105
rect 3020 65 3070 80
rect 3020 -1105 3035 65
rect 3055 -1105 3070 65
rect 3020 -1120 3070 -1105
rect 3120 65 3170 80
rect 3120 -1105 3135 65
rect 3155 -1105 3170 65
rect 3120 -1120 3170 -1105
rect 3220 65 3270 80
rect 3220 -1105 3235 65
rect 3255 -1105 3270 65
rect 3220 -1120 3270 -1105
rect 3320 65 3370 80
rect 3320 -1105 3335 65
rect 3355 -1105 3370 65
rect 3320 -1120 3370 -1105
rect 3420 65 3470 80
rect 3420 -1105 3435 65
rect 3455 -1105 3470 65
rect 3420 -1120 3470 -1105
rect 3520 65 3570 80
rect 3520 -1105 3535 65
rect 3555 -1105 3570 65
rect 3520 -1120 3570 -1105
rect 3620 65 3670 80
rect 3620 -1105 3635 65
rect 3655 -1105 3670 65
rect 3620 -1120 3670 -1105
rect 3720 65 3770 80
rect 3720 -1105 3735 65
rect 3755 -1105 3770 65
rect 3720 -1120 3770 -1105
rect 3820 65 3870 80
rect 3820 -1105 3835 65
rect 3855 -1105 3870 65
rect 3820 -1120 3870 -1105
rect 3920 65 3970 80
rect 3920 -1105 3935 65
rect 3955 -1105 3970 65
rect 3920 -1120 3970 -1105
rect 4020 65 4070 80
rect 4020 -1105 4035 65
rect 4055 -1105 4070 65
rect 4020 -1120 4070 -1105
<< ndiffc >>
rect 810 -2435 830 -1270
rect 910 -2435 930 -1270
rect 1040 -2440 1060 -1270
rect 1140 -2440 1160 -1270
rect 1240 -2440 1260 -1270
rect 1340 -2440 1360 -1270
rect 1440 -2440 1460 -1270
rect 1540 -2440 1560 -1270
rect 1640 -2440 1660 -1270
rect 1740 -2440 1760 -1270
rect 1840 -2440 1860 -1270
rect 1940 -2440 1960 -1270
rect 2040 -2440 2060 -1270
rect 2140 -2440 2160 -1270
rect 2240 -2440 2260 -1270
rect 2340 -2440 2360 -1270
rect 2440 -2440 2460 -1270
rect 2635 -2440 2655 -1270
rect 2735 -2440 2755 -1270
rect 2835 -2440 2855 -1270
rect 2935 -2440 2955 -1270
rect 3035 -2440 3055 -1270
rect 3135 -2440 3155 -1270
rect 3235 -2440 3255 -1270
rect 3335 -2440 3355 -1270
rect 3435 -2440 3455 -1270
rect 3535 -2440 3555 -1270
rect 3635 -2440 3655 -1270
rect 3735 -2440 3755 -1270
rect 3835 -2440 3855 -1270
rect 3935 -2440 3955 -1270
rect 4035 -2440 4055 -1270
<< pdiffc >>
rect 620 65 890 85
rect 620 -35 890 -15
rect 620 -135 890 -115
rect 620 -235 890 -215
rect 620 -335 890 -315
rect 620 -435 890 -415
rect 620 -535 890 -515
rect 620 -635 890 -615
rect 620 -735 890 -715
rect 620 -835 890 -815
rect 620 -935 890 -915
rect 1040 -1040 1060 130
rect 1140 -1040 1160 130
rect 1240 -1040 1260 130
rect 1340 -1040 1360 130
rect 1440 -1040 1460 130
rect 1540 -1040 1560 130
rect 1640 -1040 1660 130
rect 1740 -1040 1760 130
rect 1840 -1040 1860 130
rect 1940 -1040 1960 130
rect 2040 -1040 2060 130
rect 2140 -1040 2160 130
rect 2240 -1040 2260 130
rect 2340 -1040 2360 130
rect 2440 -1040 2460 130
rect 2635 -1105 2655 65
rect 2735 -1105 2755 65
rect 2835 -1105 2855 65
rect 2935 -1105 2955 65
rect 3035 -1105 3055 65
rect 3135 -1105 3155 65
rect 3235 -1105 3255 65
rect 3335 -1105 3355 65
rect 3435 -1105 3455 65
rect 3535 -1105 3555 65
rect 3635 -1105 3655 65
rect 3735 -1105 3755 65
rect 3835 -1105 3855 65
rect 3935 -1105 3955 65
rect 4035 -1105 4055 65
<< psubdiff >>
rect 975 -1270 1025 -1255
rect 975 -2440 990 -1270
rect 1010 -2440 1025 -1270
rect 975 -2455 1025 -2440
rect 2470 -1270 2520 -1255
rect 2470 -2440 2485 -1270
rect 2505 -2440 2520 -1270
rect 2470 -2455 2520 -2440
rect 2575 -1270 2625 -1255
rect 2575 -2440 2590 -1270
rect 2610 -2440 2625 -1270
rect 2575 -2455 2625 -2440
rect 4070 -1270 4120 -1255
rect 4070 -2440 4085 -1270
rect 4105 -2440 4120 -1270
rect 4070 -2455 4120 -2440
<< nsubdiff >>
rect 605 130 905 145
rect 605 110 620 130
rect 890 110 905 130
rect 605 95 905 110
rect 975 130 1025 145
rect 605 -965 905 -950
rect 605 -985 620 -965
rect 890 -985 905 -965
rect 605 -1000 905 -985
rect 975 -1040 990 130
rect 1010 -1040 1025 130
rect 975 -1055 1025 -1040
rect 2470 130 2520 145
rect 2470 -1040 2485 130
rect 2505 -1040 2520 130
rect 2470 -1055 2520 -1040
rect 2575 65 2625 80
rect 2575 -1105 2590 65
rect 2610 -1105 2625 65
rect 2575 -1120 2625 -1105
rect 4070 65 4120 80
rect 4070 -1105 4085 65
rect 4105 -1105 4120 65
rect 4070 -1120 4120 -1105
<< psubdiffcont >>
rect 990 -2440 1010 -1270
rect 2485 -2440 2505 -1270
rect 2590 -2440 2610 -1270
rect 4085 -2440 4105 -1270
<< nsubdiffcont >>
rect 620 110 890 130
rect 620 -985 890 -965
rect 990 -1040 1010 130
rect 2485 -1040 2505 130
rect 2590 -1105 2610 65
rect 4085 -1105 4105 65
<< poly >>
rect 1175 190 1225 200
rect 1175 170 1190 190
rect 1210 170 1225 190
rect 1075 145 1125 160
rect 1175 145 1225 170
rect 1275 190 1325 200
rect 1275 170 1290 190
rect 1310 170 1325 190
rect 1275 145 1325 170
rect 1375 190 1425 200
rect 1375 170 1390 190
rect 1410 170 1425 190
rect 1375 145 1425 170
rect 1475 190 1525 200
rect 1475 170 1490 190
rect 1510 170 1525 190
rect 1475 145 1525 170
rect 1575 190 1625 200
rect 1575 170 1590 190
rect 1610 170 1625 190
rect 1575 145 1625 170
rect 1675 190 1725 200
rect 1675 170 1690 190
rect 1710 170 1725 190
rect 1675 145 1725 170
rect 1775 190 1825 200
rect 1775 170 1790 190
rect 1810 170 1825 190
rect 1775 145 1825 170
rect 1875 190 1925 200
rect 1875 170 1890 190
rect 1910 170 1925 190
rect 1875 145 1925 170
rect 1975 190 2025 200
rect 1975 170 1990 190
rect 2010 170 2025 190
rect 1975 145 2025 170
rect 2075 190 2125 200
rect 2075 170 2090 190
rect 2110 170 2125 190
rect 2075 145 2125 170
rect 2175 190 2225 200
rect 2175 170 2190 190
rect 2210 170 2225 190
rect 2175 145 2225 170
rect 2275 190 2325 200
rect 2275 170 2290 190
rect 2310 170 2325 190
rect 2275 145 2325 170
rect 2375 145 2425 160
rect 920 50 960 55
rect 590 0 605 50
rect 905 45 960 50
rect 905 25 930 45
rect 950 25 960 45
rect 905 0 960 25
rect 550 -65 605 -50
rect 550 -85 560 -65
rect 580 -85 605 -65
rect 550 -100 605 -85
rect 905 -100 920 -50
rect 550 -165 605 -150
rect 550 -185 560 -165
rect 580 -185 605 -165
rect 550 -200 605 -185
rect 905 -200 920 -150
rect 550 -265 605 -250
rect 550 -285 560 -265
rect 580 -285 605 -265
rect 550 -300 605 -285
rect 905 -300 920 -250
rect 550 -365 605 -350
rect 550 -385 560 -365
rect 580 -385 605 -365
rect 550 -400 605 -385
rect 905 -400 920 -350
rect 550 -465 605 -450
rect 550 -485 560 -465
rect 580 -485 605 -465
rect 550 -500 605 -485
rect 905 -500 920 -450
rect 550 -565 605 -550
rect 550 -585 560 -565
rect 580 -585 605 -565
rect 550 -600 605 -585
rect 905 -600 920 -550
rect 550 -665 605 -650
rect 550 -685 560 -665
rect 580 -685 605 -665
rect 550 -700 605 -685
rect 905 -700 920 -650
rect 550 -775 605 -750
rect 550 -795 560 -775
rect 580 -795 605 -775
rect 550 -800 605 -795
rect 905 -800 920 -750
rect 550 -805 590 -800
rect 550 -865 605 -850
rect 550 -885 560 -865
rect 580 -885 605 -865
rect 550 -900 605 -885
rect 905 -900 920 -850
rect 2665 135 2720 145
rect 2665 115 2675 135
rect 2695 115 2720 135
rect 2665 105 2720 115
rect 2670 80 2720 105
rect 3970 135 4025 145
rect 3970 115 3995 135
rect 4015 115 4025 135
rect 3970 105 4025 115
rect 2770 80 2820 100
rect 2870 80 2920 100
rect 2970 80 3020 100
rect 3070 80 3120 100
rect 3170 80 3220 100
rect 3270 80 3320 100
rect 3370 80 3420 100
rect 3470 80 3520 100
rect 3570 80 3620 100
rect 3670 80 3720 100
rect 3770 80 3820 100
rect 3870 80 3920 100
rect 3970 80 4020 105
rect 1075 -1080 1125 -1055
rect 1175 -1075 1225 -1055
rect 1275 -1075 1325 -1055
rect 1375 -1075 1425 -1055
rect 1475 -1075 1525 -1055
rect 1575 -1075 1625 -1055
rect 1675 -1075 1725 -1055
rect 1775 -1075 1825 -1055
rect 1875 -1075 1925 -1055
rect 1975 -1075 2025 -1055
rect 2075 -1075 2125 -1055
rect 2175 -1075 2225 -1055
rect 2275 -1075 2325 -1055
rect 1070 -1090 1125 -1080
rect 1070 -1110 1080 -1090
rect 1100 -1110 1125 -1090
rect 1070 -1120 1125 -1110
rect 2375 -1080 2425 -1055
rect 2375 -1090 2430 -1080
rect 2375 -1110 2400 -1090
rect 2420 -1110 2430 -1090
rect 2375 -1120 2430 -1110
rect 2670 -1135 2720 -1120
rect 2770 -1145 2820 -1120
rect 2770 -1165 2785 -1145
rect 2805 -1165 2820 -1145
rect 2770 -1175 2820 -1165
rect 2870 -1145 2920 -1120
rect 2870 -1165 2885 -1145
rect 2905 -1165 2920 -1145
rect 2870 -1175 2920 -1165
rect 2970 -1145 3020 -1120
rect 2970 -1165 2985 -1145
rect 3005 -1165 3020 -1145
rect 2970 -1175 3020 -1165
rect 3070 -1145 3120 -1120
rect 3070 -1165 3085 -1145
rect 3105 -1165 3120 -1145
rect 3070 -1175 3120 -1165
rect 3170 -1145 3220 -1120
rect 3170 -1165 3185 -1145
rect 3205 -1165 3220 -1145
rect 3170 -1175 3220 -1165
rect 3270 -1145 3320 -1120
rect 3270 -1165 3285 -1145
rect 3305 -1165 3320 -1145
rect 3270 -1175 3320 -1165
rect 3370 -1145 3420 -1120
rect 3370 -1165 3385 -1145
rect 3405 -1165 3420 -1145
rect 3370 -1175 3420 -1165
rect 3470 -1145 3520 -1120
rect 3470 -1165 3485 -1145
rect 3505 -1165 3520 -1145
rect 3470 -1175 3520 -1165
rect 3570 -1145 3620 -1120
rect 3570 -1165 3585 -1145
rect 3605 -1165 3620 -1145
rect 3570 -1175 3620 -1165
rect 3670 -1145 3720 -1120
rect 3670 -1165 3685 -1145
rect 3705 -1165 3720 -1145
rect 3670 -1175 3720 -1165
rect 3770 -1145 3820 -1120
rect 3770 -1165 3785 -1145
rect 3805 -1165 3820 -1145
rect 3770 -1175 3820 -1165
rect 3870 -1145 3920 -1120
rect 3970 -1135 4020 -1120
rect 3870 -1165 3885 -1145
rect 3905 -1165 3920 -1145
rect 3870 -1175 3920 -1165
rect 2665 -1200 2720 -1190
rect 1175 -1210 1225 -1200
rect 1175 -1230 1190 -1210
rect 1210 -1230 1225 -1210
rect 845 -1255 895 -1240
rect 1075 -1255 1125 -1240
rect 1175 -1255 1225 -1230
rect 1275 -1210 1325 -1200
rect 1275 -1230 1290 -1210
rect 1310 -1230 1325 -1210
rect 1275 -1255 1325 -1230
rect 1375 -1210 1425 -1200
rect 1375 -1230 1390 -1210
rect 1410 -1230 1425 -1210
rect 1375 -1255 1425 -1230
rect 1475 -1210 1525 -1200
rect 1475 -1230 1490 -1210
rect 1510 -1230 1525 -1210
rect 1475 -1255 1525 -1230
rect 1575 -1210 1625 -1200
rect 1575 -1230 1590 -1210
rect 1610 -1230 1625 -1210
rect 1575 -1255 1625 -1230
rect 1675 -1210 1725 -1200
rect 1675 -1230 1690 -1210
rect 1710 -1230 1725 -1210
rect 1675 -1255 1725 -1230
rect 1775 -1210 1825 -1200
rect 1775 -1230 1790 -1210
rect 1810 -1230 1825 -1210
rect 1775 -1255 1825 -1230
rect 1875 -1210 1925 -1200
rect 1875 -1230 1890 -1210
rect 1910 -1230 1925 -1210
rect 1875 -1255 1925 -1230
rect 1975 -1210 2025 -1200
rect 1975 -1230 1990 -1210
rect 2010 -1230 2025 -1210
rect 1975 -1255 2025 -1230
rect 2075 -1210 2125 -1200
rect 2075 -1230 2090 -1210
rect 2110 -1230 2125 -1210
rect 2075 -1255 2125 -1230
rect 2175 -1210 2225 -1200
rect 2175 -1230 2190 -1210
rect 2210 -1230 2225 -1210
rect 2175 -1255 2225 -1230
rect 2275 -1210 2325 -1200
rect 2275 -1230 2290 -1210
rect 2310 -1230 2325 -1210
rect 2665 -1220 2675 -1200
rect 2695 -1220 2720 -1200
rect 2665 -1230 2720 -1220
rect 2275 -1255 2325 -1230
rect 2375 -1255 2425 -1240
rect 2670 -1255 2720 -1230
rect 3970 -1200 4025 -1190
rect 3970 -1220 3995 -1200
rect 4015 -1220 4025 -1200
rect 3970 -1230 4025 -1220
rect 2770 -1255 2820 -1235
rect 2870 -1255 2920 -1235
rect 2970 -1255 3020 -1235
rect 3070 -1255 3120 -1235
rect 3170 -1255 3220 -1235
rect 3270 -1255 3320 -1235
rect 3370 -1255 3420 -1235
rect 3470 -1255 3520 -1235
rect 3570 -1255 3620 -1235
rect 3670 -1255 3720 -1235
rect 3770 -1255 3820 -1235
rect 3870 -1255 3920 -1235
rect 3970 -1255 4020 -1230
rect 845 -2475 895 -2455
rect 845 -2495 855 -2475
rect 875 -2495 895 -2475
rect 1075 -2480 1125 -2455
rect 1175 -2475 1225 -2455
rect 1275 -2475 1325 -2455
rect 1375 -2475 1425 -2455
rect 1475 -2475 1525 -2455
rect 1575 -2475 1625 -2455
rect 1675 -2475 1725 -2455
rect 1775 -2475 1825 -2455
rect 1875 -2475 1925 -2455
rect 1975 -2475 2025 -2455
rect 2075 -2475 2125 -2455
rect 2175 -2475 2225 -2455
rect 2275 -2475 2325 -2455
rect 845 -2505 895 -2495
rect 1070 -2490 1125 -2480
rect 1070 -2510 1080 -2490
rect 1100 -2510 1125 -2490
rect 1070 -2520 1125 -2510
rect 2375 -2480 2425 -2455
rect 2670 -2470 2720 -2455
rect 2770 -2480 2820 -2455
rect 2375 -2490 2430 -2480
rect 2375 -2510 2400 -2490
rect 2420 -2510 2430 -2490
rect 2770 -2500 2785 -2480
rect 2805 -2500 2820 -2480
rect 2770 -2510 2820 -2500
rect 2870 -2480 2920 -2455
rect 2870 -2500 2885 -2480
rect 2905 -2500 2920 -2480
rect 2870 -2510 2920 -2500
rect 2970 -2480 3020 -2455
rect 2970 -2500 2985 -2480
rect 3005 -2500 3020 -2480
rect 2970 -2510 3020 -2500
rect 3070 -2480 3120 -2455
rect 3070 -2500 3085 -2480
rect 3105 -2500 3120 -2480
rect 3070 -2510 3120 -2500
rect 3170 -2480 3220 -2455
rect 3170 -2500 3185 -2480
rect 3205 -2500 3220 -2480
rect 3170 -2510 3220 -2500
rect 3270 -2480 3320 -2455
rect 3270 -2500 3285 -2480
rect 3305 -2500 3320 -2480
rect 3270 -2510 3320 -2500
rect 3370 -2480 3420 -2455
rect 3370 -2500 3385 -2480
rect 3405 -2500 3420 -2480
rect 3370 -2510 3420 -2500
rect 3470 -2480 3520 -2455
rect 3470 -2500 3485 -2480
rect 3505 -2500 3520 -2480
rect 3470 -2510 3520 -2500
rect 3570 -2480 3620 -2455
rect 3570 -2500 3585 -2480
rect 3605 -2500 3620 -2480
rect 3570 -2510 3620 -2500
rect 3670 -2480 3720 -2455
rect 3670 -2500 3685 -2480
rect 3705 -2500 3720 -2480
rect 3670 -2510 3720 -2500
rect 3770 -2480 3820 -2455
rect 3770 -2500 3785 -2480
rect 3805 -2500 3820 -2480
rect 3770 -2510 3820 -2500
rect 3870 -2480 3920 -2455
rect 3970 -2470 4020 -2455
rect 3870 -2500 3885 -2480
rect 3905 -2500 3920 -2480
rect 3870 -2510 3920 -2500
rect 2375 -2520 2430 -2510
<< polycont >>
rect 1190 170 1210 190
rect 1290 170 1310 190
rect 1390 170 1410 190
rect 1490 170 1510 190
rect 1590 170 1610 190
rect 1690 170 1710 190
rect 1790 170 1810 190
rect 1890 170 1910 190
rect 1990 170 2010 190
rect 2090 170 2110 190
rect 2190 170 2210 190
rect 2290 170 2310 190
rect 930 25 950 45
rect 560 -85 580 -65
rect 560 -185 580 -165
rect 560 -285 580 -265
rect 560 -385 580 -365
rect 560 -485 580 -465
rect 560 -585 580 -565
rect 560 -685 580 -665
rect 560 -795 580 -775
rect 560 -885 580 -865
rect 2675 115 2695 135
rect 3995 115 4015 135
rect 1080 -1110 1100 -1090
rect 2400 -1110 2420 -1090
rect 2785 -1165 2805 -1145
rect 2885 -1165 2905 -1145
rect 2985 -1165 3005 -1145
rect 3085 -1165 3105 -1145
rect 3185 -1165 3205 -1145
rect 3285 -1165 3305 -1145
rect 3385 -1165 3405 -1145
rect 3485 -1165 3505 -1145
rect 3585 -1165 3605 -1145
rect 3685 -1165 3705 -1145
rect 3785 -1165 3805 -1145
rect 3885 -1165 3905 -1145
rect 1190 -1230 1210 -1210
rect 1290 -1230 1310 -1210
rect 1390 -1230 1410 -1210
rect 1490 -1230 1510 -1210
rect 1590 -1230 1610 -1210
rect 1690 -1230 1710 -1210
rect 1790 -1230 1810 -1210
rect 1890 -1230 1910 -1210
rect 1990 -1230 2010 -1210
rect 2090 -1230 2110 -1210
rect 2190 -1230 2210 -1210
rect 2290 -1230 2310 -1210
rect 2675 -1220 2695 -1200
rect 3995 -1220 4015 -1200
rect 855 -2495 875 -2475
rect 1080 -2510 1100 -2490
rect 2400 -2510 2420 -2490
rect 2785 -2500 2805 -2480
rect 2885 -2500 2905 -2480
rect 2985 -2500 3005 -2480
rect 3085 -2500 3105 -2480
rect 3185 -2500 3205 -2480
rect 3285 -2500 3305 -2480
rect 3385 -2500 3405 -2480
rect 3485 -2500 3505 -2480
rect 3585 -2500 3605 -2480
rect 3685 -2500 3705 -2480
rect 3785 -2500 3805 -2480
rect 3885 -2500 3905 -2480
<< locali >>
rect 550 190 2320 200
rect 550 170 1190 190
rect 1210 170 1290 190
rect 1310 170 1390 190
rect 1410 170 1490 190
rect 1510 170 1590 190
rect 1610 170 1690 190
rect 1710 170 1790 190
rect 1810 170 1890 190
rect 1910 170 1990 190
rect 2010 170 2090 190
rect 2110 170 2190 190
rect 2210 170 2290 190
rect 2310 170 2320 190
rect 550 160 2320 170
rect 2725 160 3965 200
rect 550 -65 590 160
rect 610 130 900 140
rect 610 110 620 130
rect 890 110 900 130
rect 610 85 900 110
rect 610 65 620 85
rect 890 65 900 85
rect 610 55 900 65
rect 980 130 1070 140
rect 920 45 960 55
rect 920 25 930 45
rect 950 25 960 45
rect 920 15 960 25
rect 610 -15 960 -5
rect 610 -35 620 -15
rect 890 -35 960 -15
rect 610 -45 960 -35
rect 550 -85 560 -65
rect 580 -85 590 -65
rect 550 -165 590 -85
rect 610 -115 900 -105
rect 610 -135 620 -115
rect 890 -135 900 -115
rect 610 -145 900 -135
rect 550 -185 560 -165
rect 580 -185 590 -165
rect 550 -205 590 -185
rect 550 -215 900 -205
rect 550 -235 620 -215
rect 890 -235 900 -215
rect 550 -245 900 -235
rect 550 -265 590 -245
rect 550 -285 560 -265
rect 580 -285 590 -265
rect 550 -365 590 -285
rect 610 -315 900 -305
rect 610 -335 620 -315
rect 890 -335 900 -315
rect 610 -345 900 -335
rect 550 -385 560 -365
rect 580 -385 590 -365
rect 550 -465 590 -385
rect 920 -405 960 -45
rect 610 -415 960 -405
rect 610 -435 620 -415
rect 890 -435 960 -415
rect 610 -445 960 -435
rect 550 -485 560 -465
rect 580 -485 590 -465
rect 550 -565 590 -485
rect 610 -515 900 -505
rect 610 -535 620 -515
rect 890 -535 900 -515
rect 610 -545 900 -535
rect 550 -585 560 -565
rect 580 -585 590 -565
rect 550 -605 590 -585
rect 550 -615 900 -605
rect 550 -635 620 -615
rect 890 -635 900 -615
rect 550 -645 900 -635
rect 550 -665 590 -645
rect 550 -685 560 -665
rect 580 -685 590 -665
rect 550 -775 590 -685
rect 610 -715 900 -705
rect 610 -735 620 -715
rect 890 -735 900 -715
rect 610 -745 900 -735
rect 550 -795 560 -775
rect 580 -795 590 -775
rect 550 -805 590 -795
rect 920 -805 960 -445
rect 610 -815 960 -805
rect 610 -835 620 -815
rect 890 -835 960 -815
rect 610 -845 960 -835
rect 550 -865 590 -855
rect 550 -885 560 -865
rect 580 -885 590 -865
rect 550 -895 590 -885
rect 610 -915 900 -905
rect 610 -935 620 -915
rect 890 -935 900 -915
rect 610 -965 900 -935
rect 610 -985 620 -965
rect 890 -985 900 -965
rect 610 -995 900 -985
rect 920 -1200 960 -845
rect 980 -1040 990 130
rect 1010 -1040 1040 130
rect 1060 -1040 1070 130
rect 980 -1050 1070 -1040
rect 1130 130 1170 140
rect 1130 -1040 1140 130
rect 1160 -1040 1170 130
rect 1070 -1090 1110 -1080
rect 1070 -1110 1080 -1090
rect 1100 -1110 1110 -1090
rect 1070 -1120 1110 -1110
rect 800 -1240 960 -1200
rect 1130 -1200 1170 -1040
rect 1230 130 1270 140
rect 1230 -1040 1240 130
rect 1260 -1040 1270 130
rect 1230 -1050 1270 -1040
rect 1330 130 1370 140
rect 1330 -1040 1340 130
rect 1360 -1040 1370 130
rect 1330 -1050 1370 -1040
rect 1430 130 1470 140
rect 1430 -1040 1440 130
rect 1460 -1040 1470 130
rect 1430 -1050 1470 -1040
rect 1530 130 1570 140
rect 1530 -1040 1540 130
rect 1560 -1040 1570 130
rect 1530 -1050 1570 -1040
rect 1630 130 1670 140
rect 1630 -1040 1640 130
rect 1660 -1040 1670 130
rect 1630 -1050 1670 -1040
rect 1730 130 1770 140
rect 1730 -1040 1740 130
rect 1760 -1040 1770 130
rect 1730 -1200 1770 -1040
rect 1830 130 1870 140
rect 1830 -1040 1840 130
rect 1860 -1040 1870 130
rect 1830 -1050 1870 -1040
rect 1930 130 1970 140
rect 1930 -1040 1940 130
rect 1960 -1040 1970 130
rect 1930 -1050 1970 -1040
rect 2030 130 2070 140
rect 2030 -1040 2040 130
rect 2060 -1040 2070 130
rect 2030 -1050 2070 -1040
rect 2130 130 2170 140
rect 2130 -1040 2140 130
rect 2160 -1040 2170 130
rect 2130 -1050 2170 -1040
rect 2230 130 2270 140
rect 2230 -1040 2240 130
rect 2260 -1040 2270 130
rect 2230 -1050 2270 -1040
rect 2330 130 2370 140
rect 2330 -1040 2340 130
rect 2360 -1040 2370 130
rect 2330 -1200 2370 -1040
rect 2430 130 2515 140
rect 2430 -1040 2440 130
rect 2460 -1040 2485 130
rect 2505 -1040 2515 130
rect 2665 135 2705 145
rect 2665 115 2675 135
rect 2695 115 2705 135
rect 2665 105 2705 115
rect 2430 -1050 2515 -1040
rect 2580 65 2665 75
rect 2390 -1090 2430 -1080
rect 2390 -1110 2400 -1090
rect 2420 -1110 2430 -1090
rect 2390 -1120 2430 -1110
rect 2580 -1105 2590 65
rect 2610 -1105 2635 65
rect 2655 -1105 2665 65
rect 2580 -1115 2665 -1105
rect 2725 65 2765 160
rect 2725 -1105 2735 65
rect 2755 -1105 2765 65
rect 2725 -1135 2765 -1105
rect 2825 100 3865 140
rect 2825 65 2865 100
rect 2825 -1105 2835 65
rect 2855 -1105 2865 65
rect 2825 -1115 2865 -1105
rect 2925 65 2965 75
rect 2925 -1105 2935 65
rect 2955 -1105 2965 65
rect 2925 -1135 2965 -1105
rect 3025 65 3065 100
rect 3025 -1105 3035 65
rect 3055 -1105 3065 65
rect 3025 -1115 3065 -1105
rect 3125 65 3165 75
rect 3125 -1105 3135 65
rect 3155 -1105 3165 65
rect 3125 -1135 3165 -1105
rect 3225 65 3265 100
rect 3225 -1105 3235 65
rect 3255 -1105 3265 65
rect 3225 -1115 3265 -1105
rect 3325 65 3365 75
rect 3325 -1105 3335 65
rect 3355 -1105 3365 65
rect 3325 -1115 3365 -1105
rect 3425 65 3465 100
rect 3425 -1105 3435 65
rect 3455 -1105 3465 65
rect 3425 -1115 3465 -1105
rect 3525 65 3565 75
rect 3525 -1105 3535 65
rect 3555 -1105 3565 65
rect 3525 -1135 3565 -1105
rect 3625 65 3665 100
rect 3625 -1105 3635 65
rect 3655 -1105 3665 65
rect 3625 -1115 3665 -1105
rect 3725 65 3765 75
rect 3725 -1105 3735 65
rect 3755 -1105 3765 65
rect 3725 -1135 3765 -1105
rect 3825 65 3865 100
rect 3825 -1105 3835 65
rect 3855 -1105 3865 65
rect 3825 -1115 3865 -1105
rect 3925 65 3965 160
rect 3985 135 4025 145
rect 3985 115 3995 135
rect 4015 115 4025 135
rect 3985 105 4025 115
rect 3925 -1105 3935 65
rect 3955 -1105 3965 65
rect 3925 -1135 3965 -1105
rect 4025 65 4115 75
rect 4025 -1105 4035 65
rect 4055 -1105 4085 65
rect 4105 -1105 4115 65
rect 4025 -1115 4115 -1105
rect 2725 -1145 2815 -1135
rect 2725 -1165 2785 -1145
rect 2805 -1165 2815 -1145
rect 2725 -1175 2815 -1165
rect 2875 -1145 3815 -1135
rect 2875 -1165 2885 -1145
rect 2905 -1165 2985 -1145
rect 3005 -1165 3085 -1145
rect 3105 -1165 3185 -1145
rect 3205 -1165 3285 -1145
rect 3305 -1165 3385 -1145
rect 3405 -1165 3485 -1145
rect 3505 -1165 3585 -1145
rect 3605 -1165 3685 -1145
rect 3705 -1165 3785 -1145
rect 3805 -1165 3815 -1145
rect 2875 -1175 3815 -1165
rect 3875 -1145 3965 -1135
rect 3875 -1165 3885 -1145
rect 3905 -1165 3965 -1145
rect 3875 -1175 3965 -1165
rect 1130 -1210 1220 -1200
rect 1130 -1230 1190 -1210
rect 1210 -1230 1220 -1210
rect 1130 -1240 1220 -1230
rect 1280 -1210 2220 -1200
rect 1280 -1230 1290 -1210
rect 1310 -1230 1390 -1210
rect 1410 -1230 1490 -1210
rect 1510 -1230 1590 -1210
rect 1610 -1230 1690 -1210
rect 1710 -1230 1790 -1210
rect 1810 -1230 1890 -1210
rect 1910 -1230 1990 -1210
rect 2010 -1230 2090 -1210
rect 2110 -1230 2190 -1210
rect 2210 -1230 2220 -1210
rect 1280 -1240 2220 -1230
rect 2280 -1210 2370 -1200
rect 2280 -1230 2290 -1210
rect 2310 -1230 2370 -1210
rect 2665 -1200 2705 -1190
rect 2665 -1220 2675 -1200
rect 2695 -1220 2705 -1200
rect 2665 -1230 2705 -1220
rect 2280 -1240 2370 -1230
rect 800 -1270 840 -1240
rect 800 -2435 810 -1270
rect 830 -2435 840 -1270
rect 800 -2465 840 -2435
rect 900 -1270 940 -1260
rect 900 -2435 910 -1270
rect 930 -2435 940 -1270
rect 900 -2450 940 -2435
rect 980 -1270 1070 -1260
rect 980 -2440 990 -1270
rect 1010 -2440 1040 -1270
rect 1060 -2440 1070 -1270
rect 980 -2450 1070 -2440
rect 1130 -1270 1170 -1240
rect 1130 -2440 1140 -1270
rect 1160 -2440 1170 -1270
rect 800 -2475 885 -2465
rect 800 -2495 855 -2475
rect 875 -2495 885 -2475
rect 800 -2505 885 -2495
rect 1070 -2490 1110 -2480
rect 800 -2595 845 -2505
rect 1070 -2510 1080 -2490
rect 1100 -2510 1110 -2490
rect 1070 -2520 1110 -2510
rect 1130 -2535 1170 -2440
rect 1230 -1270 1270 -1260
rect 1230 -2440 1240 -1270
rect 1260 -2440 1270 -1270
rect 1230 -2475 1270 -2440
rect 1330 -1270 1370 -1240
rect 1330 -2440 1340 -1270
rect 1360 -2440 1370 -1270
rect 1330 -2450 1370 -2440
rect 1430 -1270 1470 -1260
rect 1430 -2440 1440 -1270
rect 1460 -2440 1470 -1270
rect 1430 -2475 1470 -2440
rect 1530 -1270 1570 -1240
rect 1530 -2440 1540 -1270
rect 1560 -2440 1570 -1270
rect 1530 -2450 1570 -2440
rect 1630 -1270 1670 -1260
rect 1630 -2440 1640 -1270
rect 1660 -2440 1670 -1270
rect 1630 -2475 1670 -2440
rect 1730 -1270 1770 -1260
rect 1730 -2440 1740 -1270
rect 1760 -2440 1770 -1270
rect 1730 -2450 1770 -2440
rect 1830 -1270 1870 -1260
rect 1830 -2440 1840 -1270
rect 1860 -2440 1870 -1270
rect 1830 -2475 1870 -2440
rect 1930 -1270 1970 -1240
rect 1930 -2440 1940 -1270
rect 1960 -2440 1970 -1270
rect 1930 -2450 1970 -2440
rect 2030 -1270 2070 -1260
rect 2030 -2440 2040 -1270
rect 2060 -2440 2070 -1270
rect 2030 -2475 2070 -2440
rect 2130 -1270 2170 -1240
rect 2130 -2440 2140 -1270
rect 2160 -2440 2170 -1270
rect 2130 -2450 2170 -2440
rect 2230 -1270 2270 -1260
rect 2230 -2440 2240 -1270
rect 2260 -2440 2270 -1270
rect 2230 -2475 2270 -2440
rect 1230 -2515 2270 -2475
rect 2330 -1270 2370 -1240
rect 2330 -2440 2340 -1270
rect 2360 -2440 2370 -1270
rect 2330 -2535 2370 -2440
rect 2430 -1270 2515 -1260
rect 2430 -2440 2440 -1270
rect 2460 -2440 2485 -1270
rect 2505 -2440 2515 -1270
rect 2430 -2450 2515 -2440
rect 2580 -1270 2665 -1260
rect 2580 -2440 2590 -1270
rect 2610 -2440 2635 -1270
rect 2655 -2440 2665 -1270
rect 2580 -2450 2665 -2440
rect 2725 -1270 2765 -1175
rect 2725 -2440 2735 -1270
rect 2755 -2440 2765 -1270
rect 2725 -2450 2765 -2440
rect 2825 -1270 2865 -1260
rect 2825 -2440 2835 -1270
rect 2855 -2440 2865 -1270
rect 2825 -2450 2865 -2440
rect 2925 -1270 2965 -1260
rect 2925 -2440 2935 -1270
rect 2955 -2440 2965 -1270
rect 2925 -2450 2965 -2440
rect 3025 -1270 3065 -1260
rect 3025 -2440 3035 -1270
rect 3055 -2440 3065 -1270
rect 3025 -2450 3065 -2440
rect 3125 -1270 3165 -1260
rect 3125 -2440 3135 -1270
rect 3155 -2440 3165 -1270
rect 3125 -2450 3165 -2440
rect 3225 -1270 3265 -1260
rect 3225 -2440 3235 -1270
rect 3255 -2440 3265 -1270
rect 3225 -2450 3265 -2440
rect 3325 -1270 3365 -1175
rect 3325 -2440 3335 -1270
rect 3355 -2440 3365 -1270
rect 3325 -2450 3365 -2440
rect 3425 -1270 3465 -1260
rect 3425 -2440 3435 -1270
rect 3455 -2440 3465 -1270
rect 3425 -2450 3465 -2440
rect 3525 -1270 3565 -1260
rect 3525 -2440 3535 -1270
rect 3555 -2440 3565 -1270
rect 3525 -2450 3565 -2440
rect 3625 -1270 3665 -1260
rect 3625 -2440 3635 -1270
rect 3655 -2440 3665 -1270
rect 3625 -2450 3665 -2440
rect 3725 -1270 3765 -1260
rect 3725 -2440 3735 -1270
rect 3755 -2440 3765 -1270
rect 3725 -2450 3765 -2440
rect 3825 -1270 3865 -1260
rect 3825 -2440 3835 -1270
rect 3855 -2440 3865 -1270
rect 3825 -2450 3865 -2440
rect 3925 -1270 3965 -1175
rect 3985 -1200 4025 -1190
rect 3985 -1220 3995 -1200
rect 4015 -1220 4025 -1200
rect 3985 -1230 4025 -1220
rect 3925 -2440 3935 -1270
rect 3955 -2440 3965 -1270
rect 3925 -2450 3965 -2440
rect 4025 -1270 4115 -1260
rect 4025 -2440 4035 -1270
rect 4055 -2440 4085 -1270
rect 4105 -2440 4115 -1270
rect 4025 -2450 4115 -2440
rect 2775 -2480 3915 -2470
rect 2390 -2490 2430 -2480
rect 2390 -2510 2400 -2490
rect 2420 -2510 2430 -2490
rect 2390 -2520 2430 -2510
rect 2775 -2500 2785 -2480
rect 2805 -2500 2885 -2480
rect 2905 -2500 2985 -2480
rect 3005 -2500 3085 -2480
rect 3105 -2500 3185 -2480
rect 3205 -2500 3285 -2480
rect 3305 -2500 3385 -2480
rect 3405 -2500 3485 -2480
rect 3505 -2500 3585 -2480
rect 3605 -2500 3685 -2480
rect 3705 -2500 3785 -2480
rect 3805 -2500 3885 -2480
rect 3905 -2500 3915 -2480
rect 2775 -2510 3915 -2500
rect 1130 -2575 2370 -2535
rect 2775 -2595 2820 -2510
rect 800 -2635 2820 -2595
<< viali >>
rect 620 110 890 130
rect 620 65 890 85
rect 930 25 950 45
rect 620 -135 890 -115
rect 620 -335 890 -315
rect 620 -535 890 -515
rect 620 -735 890 -715
rect 560 -885 580 -865
rect 620 -935 890 -915
rect 620 -985 890 -965
rect 990 -1040 1010 130
rect 1040 -1040 1060 130
rect 1080 -1110 1100 -1090
rect 1240 -1040 1260 130
rect 2240 -1040 2260 130
rect 2440 -1040 2460 130
rect 2485 -1040 2505 130
rect 2675 115 2695 135
rect 2400 -1110 2420 -1090
rect 2590 -1105 2610 65
rect 2635 -1105 2655 65
rect 3335 -1105 3355 65
rect 3995 115 4015 135
rect 4035 -1105 4055 65
rect 4085 -1105 4105 65
rect 2675 -1220 2695 -1200
rect 910 -2435 930 -1270
rect 990 -2440 1010 -1270
rect 1040 -2440 1060 -1270
rect 1080 -2510 1100 -2490
rect 1740 -2440 1760 -1270
rect 2440 -2440 2460 -1270
rect 2485 -2440 2505 -1270
rect 2590 -2440 2610 -1270
rect 2635 -2440 2655 -1270
rect 2835 -2440 2855 -1270
rect 3835 -2440 3855 -1270
rect 3995 -1220 4015 -1200
rect 4035 -2440 4055 -1270
rect 4085 -2440 4105 -1270
rect 2400 -2510 2420 -2490
<< metal1 >>
rect 610 130 2515 140
rect 610 110 620 130
rect 890 110 990 130
rect 610 85 990 110
rect 610 65 620 85
rect 890 65 990 85
rect 610 45 990 65
rect 610 25 930 45
rect 950 25 990 45
rect 610 -115 990 25
rect 610 -135 620 -115
rect 890 -135 990 -115
rect 610 -315 990 -135
rect 610 -335 620 -315
rect 890 -335 990 -315
rect 610 -515 990 -335
rect 610 -535 620 -515
rect 890 -535 990 -515
rect 610 -715 990 -535
rect 610 -735 620 -715
rect 890 -735 990 -715
rect 610 -855 990 -735
rect 550 -865 990 -855
rect 550 -885 560 -865
rect 580 -885 990 -865
rect 550 -895 990 -885
rect 610 -915 990 -895
rect 610 -935 620 -915
rect 890 -935 990 -915
rect 610 -965 990 -935
rect 610 -985 620 -965
rect 890 -985 990 -965
rect 610 -995 990 -985
rect 980 -1040 990 -995
rect 1010 -1040 1040 130
rect 1060 -1040 1240 130
rect 1260 -1040 2240 130
rect 2260 -1040 2440 130
rect 2460 -1040 2485 130
rect 2505 75 2515 130
rect 2665 135 2720 145
rect 2665 115 2675 135
rect 2695 115 2720 135
rect 2665 105 2720 115
rect 2670 75 2720 105
rect 3970 135 4025 145
rect 3970 115 3995 135
rect 4015 115 4025 135
rect 3970 105 4025 115
rect 3970 75 4020 105
rect 2505 65 4115 75
rect 2505 -1040 2590 65
rect 980 -1050 2590 -1040
rect 1075 -1080 1125 -1050
rect 1070 -1090 1125 -1080
rect 1070 -1110 1080 -1090
rect 1100 -1110 1125 -1090
rect 1070 -1120 1125 -1110
rect 2375 -1080 2425 -1050
rect 2375 -1090 2430 -1080
rect 2375 -1110 2400 -1090
rect 2420 -1110 2430 -1090
rect 2375 -1120 2430 -1110
rect 2580 -1105 2590 -1050
rect 2610 -1105 2635 65
rect 2655 -1105 3335 65
rect 3355 -1105 4035 65
rect 4055 -1105 4085 65
rect 4105 -1105 4115 65
rect 2580 -1115 4115 -1105
rect 2665 -1200 2720 -1190
rect 2665 -1220 2675 -1200
rect 2695 -1220 2720 -1200
rect 2665 -1230 2720 -1220
rect 2670 -1260 2720 -1230
rect 3970 -1200 4025 -1190
rect 3970 -1220 3995 -1200
rect 4015 -1220 4025 -1200
rect 3970 -1230 4025 -1220
rect 3970 -1260 4020 -1230
rect 900 -1270 4115 -1260
rect 900 -2435 910 -1270
rect 930 -2435 990 -1270
rect 900 -2440 990 -2435
rect 1010 -2440 1040 -1270
rect 1060 -2440 1740 -1270
rect 1760 -2440 2440 -1270
rect 2460 -2440 2485 -1270
rect 2505 -2440 2590 -1270
rect 2610 -2440 2635 -1270
rect 2655 -2440 2835 -1270
rect 2855 -2440 3835 -1270
rect 3855 -2440 4035 -1270
rect 4055 -2440 4085 -1270
rect 4105 -2440 4115 -1270
rect 900 -2445 4115 -2440
rect 980 -2450 4115 -2445
rect 1075 -2480 1125 -2450
rect 1070 -2490 1125 -2480
rect 1070 -2510 1080 -2490
rect 1100 -2510 1125 -2490
rect 1070 -2520 1125 -2510
rect 2375 -2480 2425 -2450
rect 2375 -2490 2430 -2480
rect 2375 -2510 2400 -2490
rect 2420 -2510 2430 -2490
rect 2375 -2520 2430 -2510
<< labels >>
rlabel locali 550 -785 550 -785 7 VBP
port 3 w
rlabel metal1 610 120 610 120 7 VP
port 1 w
rlabel locali 3965 -1230 3965 -1230 3 VCP
port 6 e
rlabel metal1 920 -1260 920 -1260 1 VN
port 2 n
rlabel locali 800 -2485 800 -2485 7 VBN
port 4 w
rlabel locali 1130 -2555 1130 -2555 7 VCN
port 5 w
<< end >>
