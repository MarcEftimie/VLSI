magic
tech sky130A
timestamp 1697332078
<< nwell >>
rect 550 -1180 4140 205
<< nmos >>
rect 845 -2555 895 -1355
rect 1075 -2555 1125 -1355
rect 1175 -2555 1225 -1355
rect 1275 -2555 1325 -1355
rect 1375 -2555 1425 -1355
rect 1475 -2555 1525 -1355
rect 1575 -2555 1625 -1355
rect 1675 -2555 1725 -1355
rect 1775 -2555 1825 -1355
rect 1875 -2555 1925 -1355
rect 1975 -2555 2025 -1355
rect 2075 -2555 2125 -1355
rect 2175 -2555 2225 -1355
rect 2275 -2555 2325 -1355
rect 2375 -2555 2425 -1355
rect 2670 -2555 2720 -1355
rect 2770 -2555 2820 -1355
rect 2870 -2555 2920 -1355
rect 2970 -2555 3020 -1355
rect 3070 -2555 3120 -1355
rect 3170 -2555 3220 -1355
rect 3270 -2555 3320 -1355
rect 3370 -2555 3420 -1355
rect 3470 -2555 3520 -1355
rect 3570 -2555 3620 -1355
rect 3670 -2555 3720 -1355
rect 3770 -2555 3820 -1355
rect 3870 -2555 3920 -1355
rect 3970 -2555 4020 -1355
<< pmos >>
rect 605 40 905 90
rect 605 -60 905 -10
rect 605 -160 905 -110
rect 605 -260 905 -210
rect 605 -360 905 -310
rect 605 -460 905 -410
rect 605 -560 905 -510
rect 605 -660 905 -610
rect 605 -760 905 -710
rect 605 -860 905 -810
rect 1075 -1055 1125 145
rect 1175 -1055 1225 145
rect 1275 -1055 1325 145
rect 1375 -1055 1425 145
rect 1475 -1055 1525 145
rect 1575 -1055 1625 145
rect 1675 -1055 1725 145
rect 1775 -1055 1825 145
rect 1875 -1055 1925 145
rect 1975 -1055 2025 145
rect 2075 -1055 2125 145
rect 2175 -1055 2225 145
rect 2275 -1055 2325 145
rect 2375 -1055 2425 145
rect 2670 -1120 2720 80
rect 2770 -1120 2820 80
rect 2870 -1120 2920 80
rect 2970 -1120 3020 80
rect 3070 -1120 3120 80
rect 3170 -1120 3220 80
rect 3270 -1120 3320 80
rect 3370 -1120 3420 80
rect 3470 -1120 3520 80
rect 3570 -1120 3620 80
rect 3670 -1120 3720 80
rect 3770 -1120 3820 80
rect 3870 -1120 3920 80
rect 3970 -1120 4020 80
<< ndiff >>
rect 795 -1370 845 -1355
rect 795 -2535 810 -1370
rect 830 -2535 845 -1370
rect 795 -2555 845 -2535
rect 895 -1370 945 -1355
rect 895 -2535 910 -1370
rect 930 -2535 945 -1370
rect 895 -2555 945 -2535
rect 1025 -1370 1075 -1355
rect 1025 -2540 1040 -1370
rect 1060 -2540 1075 -1370
rect 1025 -2555 1075 -2540
rect 1125 -1370 1175 -1355
rect 1125 -2540 1140 -1370
rect 1160 -2540 1175 -1370
rect 1125 -2555 1175 -2540
rect 1225 -1370 1275 -1355
rect 1225 -2540 1240 -1370
rect 1260 -2540 1275 -1370
rect 1225 -2555 1275 -2540
rect 1325 -1370 1375 -1355
rect 1325 -2540 1340 -1370
rect 1360 -2540 1375 -1370
rect 1325 -2555 1375 -2540
rect 1425 -1370 1475 -1355
rect 1425 -2540 1440 -1370
rect 1460 -2540 1475 -1370
rect 1425 -2555 1475 -2540
rect 1525 -1370 1575 -1355
rect 1525 -2540 1540 -1370
rect 1560 -2540 1575 -1370
rect 1525 -2555 1575 -2540
rect 1625 -1370 1675 -1355
rect 1625 -2540 1640 -1370
rect 1660 -2540 1675 -1370
rect 1625 -2555 1675 -2540
rect 1725 -1370 1775 -1355
rect 1725 -2540 1740 -1370
rect 1760 -2540 1775 -1370
rect 1725 -2555 1775 -2540
rect 1825 -1370 1875 -1355
rect 1825 -2540 1840 -1370
rect 1860 -2540 1875 -1370
rect 1825 -2555 1875 -2540
rect 1925 -1370 1975 -1355
rect 1925 -2540 1940 -1370
rect 1960 -2540 1975 -1370
rect 1925 -2555 1975 -2540
rect 2025 -1370 2075 -1355
rect 2025 -2540 2040 -1370
rect 2060 -2540 2075 -1370
rect 2025 -2555 2075 -2540
rect 2125 -1370 2175 -1355
rect 2125 -2540 2140 -1370
rect 2160 -2540 2175 -1370
rect 2125 -2555 2175 -2540
rect 2225 -1370 2275 -1355
rect 2225 -2540 2240 -1370
rect 2260 -2540 2275 -1370
rect 2225 -2555 2275 -2540
rect 2325 -1370 2375 -1355
rect 2325 -2540 2340 -1370
rect 2360 -2540 2375 -1370
rect 2325 -2555 2375 -2540
rect 2425 -1370 2470 -1355
rect 2425 -2540 2440 -1370
rect 2460 -2540 2470 -1370
rect 2425 -2555 2470 -2540
rect 2625 -1370 2670 -1355
rect 2625 -2540 2635 -1370
rect 2655 -2540 2670 -1370
rect 2625 -2555 2670 -2540
rect 2720 -1370 2770 -1355
rect 2720 -2540 2735 -1370
rect 2755 -2540 2770 -1370
rect 2720 -2555 2770 -2540
rect 2820 -1370 2870 -1355
rect 2820 -2540 2835 -1370
rect 2855 -2540 2870 -1370
rect 2820 -2555 2870 -2540
rect 2920 -1370 2970 -1355
rect 2920 -2540 2935 -1370
rect 2955 -2540 2970 -1370
rect 2920 -2555 2970 -2540
rect 3020 -1370 3070 -1355
rect 3020 -2540 3035 -1370
rect 3055 -2540 3070 -1370
rect 3020 -2555 3070 -2540
rect 3120 -1370 3170 -1355
rect 3120 -2540 3135 -1370
rect 3155 -2540 3170 -1370
rect 3120 -2555 3170 -2540
rect 3220 -1370 3270 -1355
rect 3220 -2540 3235 -1370
rect 3255 -2540 3270 -1370
rect 3220 -2555 3270 -2540
rect 3320 -1370 3370 -1355
rect 3320 -2540 3335 -1370
rect 3355 -2540 3370 -1370
rect 3320 -2555 3370 -2540
rect 3420 -1370 3470 -1355
rect 3420 -2540 3435 -1370
rect 3455 -2540 3470 -1370
rect 3420 -2555 3470 -2540
rect 3520 -1370 3570 -1355
rect 3520 -2540 3535 -1370
rect 3555 -2540 3570 -1370
rect 3520 -2555 3570 -2540
rect 3620 -1370 3670 -1355
rect 3620 -2540 3635 -1370
rect 3655 -2540 3670 -1370
rect 3620 -2555 3670 -2540
rect 3720 -1370 3770 -1355
rect 3720 -2540 3735 -1370
rect 3755 -2540 3770 -1370
rect 3720 -2555 3770 -2540
rect 3820 -1370 3870 -1355
rect 3820 -2540 3835 -1370
rect 3855 -2540 3870 -1370
rect 3820 -2555 3870 -2540
rect 3920 -1370 3970 -1355
rect 3920 -2540 3935 -1370
rect 3955 -2540 3970 -1370
rect 3920 -2555 3970 -2540
rect 4020 -1370 4070 -1355
rect 4020 -2540 4035 -1370
rect 4055 -2540 4070 -1370
rect 4020 -2555 4070 -2540
<< pdiff >>
rect 605 125 905 135
rect 605 105 620 125
rect 890 105 905 125
rect 605 90 905 105
rect 1025 130 1075 145
rect 605 25 905 40
rect 605 5 620 25
rect 890 5 905 25
rect 605 -10 905 5
rect 605 -75 905 -60
rect 605 -95 620 -75
rect 890 -95 905 -75
rect 605 -110 905 -95
rect 605 -175 905 -160
rect 605 -195 620 -175
rect 890 -195 905 -175
rect 605 -210 905 -195
rect 605 -275 905 -260
rect 605 -295 620 -275
rect 890 -295 905 -275
rect 605 -310 905 -295
rect 605 -375 905 -360
rect 605 -395 620 -375
rect 890 -395 905 -375
rect 605 -410 905 -395
rect 605 -475 905 -460
rect 605 -495 620 -475
rect 890 -495 905 -475
rect 605 -510 905 -495
rect 605 -575 905 -560
rect 605 -595 620 -575
rect 890 -595 905 -575
rect 605 -610 905 -595
rect 605 -675 905 -660
rect 605 -695 620 -675
rect 890 -695 905 -675
rect 605 -710 905 -695
rect 605 -775 905 -760
rect 605 -795 620 -775
rect 890 -795 905 -775
rect 605 -810 905 -795
rect 605 -875 905 -860
rect 605 -895 620 -875
rect 890 -895 905 -875
rect 605 -910 905 -895
rect 1025 -1040 1040 130
rect 1060 -1040 1075 130
rect 1025 -1055 1075 -1040
rect 1125 130 1175 145
rect 1125 -1040 1140 130
rect 1160 -1040 1175 130
rect 1125 -1055 1175 -1040
rect 1225 130 1275 145
rect 1225 -1040 1240 130
rect 1260 -1040 1275 130
rect 1225 -1055 1275 -1040
rect 1325 130 1375 145
rect 1325 -1040 1340 130
rect 1360 -1040 1375 130
rect 1325 -1055 1375 -1040
rect 1425 130 1475 145
rect 1425 -1040 1440 130
rect 1460 -1040 1475 130
rect 1425 -1055 1475 -1040
rect 1525 130 1575 145
rect 1525 -1040 1540 130
rect 1560 -1040 1575 130
rect 1525 -1055 1575 -1040
rect 1625 130 1675 145
rect 1625 -1040 1640 130
rect 1660 -1040 1675 130
rect 1625 -1055 1675 -1040
rect 1725 130 1775 145
rect 1725 -1040 1740 130
rect 1760 -1040 1775 130
rect 1725 -1055 1775 -1040
rect 1825 130 1875 145
rect 1825 -1040 1840 130
rect 1860 -1040 1875 130
rect 1825 -1055 1875 -1040
rect 1925 130 1975 145
rect 1925 -1040 1940 130
rect 1960 -1040 1975 130
rect 1925 -1055 1975 -1040
rect 2025 130 2075 145
rect 2025 -1040 2040 130
rect 2060 -1040 2075 130
rect 2025 -1055 2075 -1040
rect 2125 130 2175 145
rect 2125 -1040 2140 130
rect 2160 -1040 2175 130
rect 2125 -1055 2175 -1040
rect 2225 130 2275 145
rect 2225 -1040 2240 130
rect 2260 -1040 2275 130
rect 2225 -1055 2275 -1040
rect 2325 130 2375 145
rect 2325 -1040 2340 130
rect 2360 -1040 2375 130
rect 2325 -1055 2375 -1040
rect 2425 130 2470 145
rect 2425 -1040 2440 130
rect 2460 -1040 2470 130
rect 2425 -1055 2470 -1040
rect 2625 65 2670 80
rect 2625 -1105 2635 65
rect 2655 -1105 2670 65
rect 2625 -1120 2670 -1105
rect 2720 65 2770 80
rect 2720 -1105 2735 65
rect 2755 -1105 2770 65
rect 2720 -1120 2770 -1105
rect 2820 65 2870 80
rect 2820 -1105 2835 65
rect 2855 -1105 2870 65
rect 2820 -1120 2870 -1105
rect 2920 65 2970 80
rect 2920 -1105 2935 65
rect 2955 -1105 2970 65
rect 2920 -1120 2970 -1105
rect 3020 65 3070 80
rect 3020 -1105 3035 65
rect 3055 -1105 3070 65
rect 3020 -1120 3070 -1105
rect 3120 65 3170 80
rect 3120 -1105 3135 65
rect 3155 -1105 3170 65
rect 3120 -1120 3170 -1105
rect 3220 65 3270 80
rect 3220 -1105 3235 65
rect 3255 -1105 3270 65
rect 3220 -1120 3270 -1105
rect 3320 65 3370 80
rect 3320 -1105 3335 65
rect 3355 -1105 3370 65
rect 3320 -1120 3370 -1105
rect 3420 65 3470 80
rect 3420 -1105 3435 65
rect 3455 -1105 3470 65
rect 3420 -1120 3470 -1105
rect 3520 65 3570 80
rect 3520 -1105 3535 65
rect 3555 -1105 3570 65
rect 3520 -1120 3570 -1105
rect 3620 65 3670 80
rect 3620 -1105 3635 65
rect 3655 -1105 3670 65
rect 3620 -1120 3670 -1105
rect 3720 65 3770 80
rect 3720 -1105 3735 65
rect 3755 -1105 3770 65
rect 3720 -1120 3770 -1105
rect 3820 65 3870 80
rect 3820 -1105 3835 65
rect 3855 -1105 3870 65
rect 3820 -1120 3870 -1105
rect 3920 65 3970 80
rect 3920 -1105 3935 65
rect 3955 -1105 3970 65
rect 3920 -1120 3970 -1105
rect 4020 65 4070 80
rect 4020 -1105 4035 65
rect 4055 -1105 4070 65
rect 4020 -1120 4070 -1105
<< ndiffc >>
rect 810 -2535 830 -1370
rect 910 -2535 930 -1370
rect 1040 -2540 1060 -1370
rect 1140 -2540 1160 -1370
rect 1240 -2540 1260 -1370
rect 1340 -2540 1360 -1370
rect 1440 -2540 1460 -1370
rect 1540 -2540 1560 -1370
rect 1640 -2540 1660 -1370
rect 1740 -2540 1760 -1370
rect 1840 -2540 1860 -1370
rect 1940 -2540 1960 -1370
rect 2040 -2540 2060 -1370
rect 2140 -2540 2160 -1370
rect 2240 -2540 2260 -1370
rect 2340 -2540 2360 -1370
rect 2440 -2540 2460 -1370
rect 2635 -2540 2655 -1370
rect 2735 -2540 2755 -1370
rect 2835 -2540 2855 -1370
rect 2935 -2540 2955 -1370
rect 3035 -2540 3055 -1370
rect 3135 -2540 3155 -1370
rect 3235 -2540 3255 -1370
rect 3335 -2540 3355 -1370
rect 3435 -2540 3455 -1370
rect 3535 -2540 3555 -1370
rect 3635 -2540 3655 -1370
rect 3735 -2540 3755 -1370
rect 3835 -2540 3855 -1370
rect 3935 -2540 3955 -1370
rect 4035 -2540 4055 -1370
<< pdiffc >>
rect 620 105 890 125
rect 620 5 890 25
rect 620 -95 890 -75
rect 620 -195 890 -175
rect 620 -295 890 -275
rect 620 -395 890 -375
rect 620 -495 890 -475
rect 620 -595 890 -575
rect 620 -695 890 -675
rect 620 -795 890 -775
rect 620 -895 890 -875
rect 1040 -1040 1060 130
rect 1140 -1040 1160 130
rect 1240 -1040 1260 130
rect 1340 -1040 1360 130
rect 1440 -1040 1460 130
rect 1540 -1040 1560 130
rect 1640 -1040 1660 130
rect 1740 -1040 1760 130
rect 1840 -1040 1860 130
rect 1940 -1040 1960 130
rect 2040 -1040 2060 130
rect 2140 -1040 2160 130
rect 2240 -1040 2260 130
rect 2340 -1040 2360 130
rect 2440 -1040 2460 130
rect 2635 -1105 2655 65
rect 2735 -1105 2755 65
rect 2835 -1105 2855 65
rect 2935 -1105 2955 65
rect 3035 -1105 3055 65
rect 3135 -1105 3155 65
rect 3235 -1105 3255 65
rect 3335 -1105 3355 65
rect 3435 -1105 3455 65
rect 3535 -1105 3555 65
rect 3635 -1105 3655 65
rect 3735 -1105 3755 65
rect 3835 -1105 3855 65
rect 3935 -1105 3955 65
rect 4035 -1105 4055 65
<< psubdiff >>
rect 975 -1370 1025 -1355
rect 975 -2540 990 -1370
rect 1010 -2540 1025 -1370
rect 975 -2555 1025 -2540
rect 2470 -1370 2520 -1355
rect 2470 -2540 2485 -1370
rect 2505 -2540 2520 -1370
rect 2470 -2555 2520 -2540
rect 2575 -1370 2625 -1355
rect 2575 -2540 2590 -1370
rect 2610 -2540 2625 -1370
rect 2575 -2555 2625 -2540
rect 4070 -1370 4120 -1355
rect 4070 -2540 4085 -1370
rect 4105 -2540 4120 -1370
rect 4070 -2555 4120 -2540
<< nsubdiff >>
rect 605 170 905 185
rect 605 150 620 170
rect 890 150 905 170
rect 605 135 905 150
rect 975 130 1025 145
rect 605 -925 905 -910
rect 605 -945 620 -925
rect 890 -945 905 -925
rect 605 -960 905 -945
rect 975 -1040 990 130
rect 1010 -1040 1025 130
rect 975 -1055 1025 -1040
rect 2470 130 2520 145
rect 2470 -1040 2485 130
rect 2505 -1040 2520 130
rect 2470 -1055 2520 -1040
rect 2575 65 2625 80
rect 2575 -1105 2590 65
rect 2610 -1105 2625 65
rect 2575 -1120 2625 -1105
rect 4070 65 4120 80
rect 4070 -1105 4085 65
rect 4105 -1105 4120 65
rect 4070 -1120 4120 -1105
<< psubdiffcont >>
rect 990 -2540 1010 -1370
rect 2485 -2540 2505 -1370
rect 2590 -2540 2610 -1370
rect 4085 -2540 4105 -1370
<< nsubdiffcont >>
rect 620 150 890 170
rect 620 -945 890 -925
rect 990 -1040 1010 130
rect 2485 -1040 2505 130
rect 2590 -1105 2610 65
rect 4085 -1105 4105 65
<< poly >>
rect 1175 190 1225 200
rect 1175 170 1190 190
rect 1210 170 1225 190
rect 1075 145 1125 160
rect 1175 145 1225 170
rect 1275 190 1325 200
rect 1275 170 1290 190
rect 1310 170 1325 190
rect 1275 145 1325 170
rect 1375 190 1425 200
rect 1375 170 1390 190
rect 1410 170 1425 190
rect 1375 145 1425 170
rect 1475 190 1525 200
rect 1475 170 1490 190
rect 1510 170 1525 190
rect 1475 145 1525 170
rect 1575 190 1625 200
rect 1575 170 1590 190
rect 1610 170 1625 190
rect 1575 145 1625 170
rect 1675 190 1725 200
rect 1675 170 1690 190
rect 1710 170 1725 190
rect 1675 145 1725 170
rect 1775 190 1825 200
rect 1775 170 1790 190
rect 1810 170 1825 190
rect 1775 145 1825 170
rect 1875 190 1925 200
rect 1875 170 1890 190
rect 1910 170 1925 190
rect 1875 145 1925 170
rect 1975 190 2025 200
rect 1975 170 1990 190
rect 2010 170 2025 190
rect 1975 145 2025 170
rect 2075 190 2125 200
rect 2075 170 2090 190
rect 2110 170 2125 190
rect 2075 145 2125 170
rect 2175 190 2225 200
rect 2175 170 2190 190
rect 2210 170 2225 190
rect 2175 145 2225 170
rect 2275 190 2325 200
rect 2275 170 2290 190
rect 2310 170 2325 190
rect 2275 145 2325 170
rect 2375 145 2425 160
rect 550 75 605 90
rect 550 55 560 75
rect 580 55 605 75
rect 550 40 605 55
rect 905 40 920 90
rect 550 -25 605 -10
rect 550 -45 560 -25
rect 580 -45 605 -25
rect 550 -60 605 -45
rect 905 -60 920 -10
rect 550 -125 605 -110
rect 550 -145 560 -125
rect 580 -145 605 -125
rect 550 -160 605 -145
rect 905 -160 920 -110
rect 550 -225 605 -210
rect 550 -245 560 -225
rect 580 -245 605 -225
rect 550 -260 605 -245
rect 905 -260 920 -210
rect 550 -325 605 -310
rect 550 -345 560 -325
rect 580 -345 605 -325
rect 550 -360 605 -345
rect 905 -360 920 -310
rect 550 -425 605 -410
rect 550 -445 560 -425
rect 580 -445 605 -425
rect 550 -460 605 -445
rect 905 -460 920 -410
rect 550 -525 605 -510
rect 550 -545 560 -525
rect 580 -545 605 -525
rect 550 -560 605 -545
rect 905 -560 920 -510
rect 550 -625 605 -610
rect 550 -645 560 -625
rect 580 -645 605 -625
rect 550 -660 605 -645
rect 905 -660 920 -610
rect 550 -735 605 -710
rect 550 -755 560 -735
rect 580 -755 605 -735
rect 550 -760 605 -755
rect 905 -760 920 -710
rect 550 -765 590 -760
rect 550 -825 605 -810
rect 550 -845 560 -825
rect 580 -845 605 -825
rect 550 -860 605 -845
rect 905 -860 920 -810
rect 2665 135 2720 145
rect 2665 115 2675 135
rect 2695 115 2720 135
rect 2665 105 2720 115
rect 2670 80 2720 105
rect 3970 135 4025 145
rect 3970 115 3995 135
rect 4015 115 4025 135
rect 3970 105 4025 115
rect 2770 80 2820 100
rect 2870 80 2920 100
rect 2970 80 3020 100
rect 3070 80 3120 100
rect 3170 80 3220 100
rect 3270 80 3320 100
rect 3370 80 3420 100
rect 3470 80 3520 100
rect 3570 80 3620 100
rect 3670 80 3720 100
rect 3770 80 3820 100
rect 3870 80 3920 100
rect 3970 80 4020 105
rect 1075 -1080 1125 -1055
rect 1175 -1075 1225 -1055
rect 1275 -1075 1325 -1055
rect 1375 -1075 1425 -1055
rect 1475 -1075 1525 -1055
rect 1575 -1075 1625 -1055
rect 1675 -1075 1725 -1055
rect 1775 -1075 1825 -1055
rect 1875 -1075 1925 -1055
rect 1975 -1075 2025 -1055
rect 2075 -1075 2125 -1055
rect 2175 -1075 2225 -1055
rect 2275 -1075 2325 -1055
rect 1070 -1090 1125 -1080
rect 1070 -1110 1080 -1090
rect 1100 -1110 1125 -1090
rect 1070 -1120 1125 -1110
rect 2375 -1080 2425 -1055
rect 2375 -1090 2430 -1080
rect 2375 -1110 2400 -1090
rect 2420 -1110 2430 -1090
rect 2375 -1120 2430 -1110
rect 2670 -1135 2720 -1120
rect 2770 -1145 2820 -1120
rect 2770 -1165 2785 -1145
rect 2805 -1165 2820 -1145
rect 2770 -1175 2820 -1165
rect 2870 -1145 2920 -1120
rect 2870 -1165 2885 -1145
rect 2905 -1165 2920 -1145
rect 2870 -1175 2920 -1165
rect 2970 -1145 3020 -1120
rect 2970 -1165 2985 -1145
rect 3005 -1165 3020 -1145
rect 2970 -1175 3020 -1165
rect 3070 -1145 3120 -1120
rect 3070 -1165 3085 -1145
rect 3105 -1165 3120 -1145
rect 3070 -1175 3120 -1165
rect 3170 -1145 3220 -1120
rect 3170 -1165 3185 -1145
rect 3205 -1165 3220 -1145
rect 3170 -1175 3220 -1165
rect 3270 -1145 3320 -1120
rect 3270 -1165 3285 -1145
rect 3305 -1165 3320 -1145
rect 3270 -1175 3320 -1165
rect 3370 -1145 3420 -1120
rect 3370 -1165 3385 -1145
rect 3405 -1165 3420 -1145
rect 3370 -1175 3420 -1165
rect 3470 -1145 3520 -1120
rect 3470 -1165 3485 -1145
rect 3505 -1165 3520 -1145
rect 3470 -1175 3520 -1165
rect 3570 -1145 3620 -1120
rect 3570 -1165 3585 -1145
rect 3605 -1165 3620 -1145
rect 3570 -1175 3620 -1165
rect 3670 -1145 3720 -1120
rect 3670 -1165 3685 -1145
rect 3705 -1165 3720 -1145
rect 3670 -1175 3720 -1165
rect 3770 -1145 3820 -1120
rect 3770 -1165 3785 -1145
rect 3805 -1165 3820 -1145
rect 3770 -1175 3820 -1165
rect 3870 -1145 3920 -1120
rect 3970 -1135 4020 -1120
rect 3870 -1165 3885 -1145
rect 3905 -1165 3920 -1145
rect 3870 -1175 3920 -1165
rect 2665 -1300 2720 -1290
rect 1175 -1310 1225 -1300
rect 1175 -1330 1190 -1310
rect 1210 -1330 1225 -1310
rect 845 -1355 895 -1340
rect 1075 -1355 1125 -1340
rect 1175 -1355 1225 -1330
rect 1275 -1310 1325 -1300
rect 1275 -1330 1290 -1310
rect 1310 -1330 1325 -1310
rect 1275 -1355 1325 -1330
rect 1375 -1310 1425 -1300
rect 1375 -1330 1390 -1310
rect 1410 -1330 1425 -1310
rect 1375 -1355 1425 -1330
rect 1475 -1310 1525 -1300
rect 1475 -1330 1490 -1310
rect 1510 -1330 1525 -1310
rect 1475 -1355 1525 -1330
rect 1575 -1310 1625 -1300
rect 1575 -1330 1590 -1310
rect 1610 -1330 1625 -1310
rect 1575 -1355 1625 -1330
rect 1675 -1310 1725 -1300
rect 1675 -1330 1690 -1310
rect 1710 -1330 1725 -1310
rect 1675 -1355 1725 -1330
rect 1775 -1310 1825 -1300
rect 1775 -1330 1790 -1310
rect 1810 -1330 1825 -1310
rect 1775 -1355 1825 -1330
rect 1875 -1310 1925 -1300
rect 1875 -1330 1890 -1310
rect 1910 -1330 1925 -1310
rect 1875 -1355 1925 -1330
rect 1975 -1310 2025 -1300
rect 1975 -1330 1990 -1310
rect 2010 -1330 2025 -1310
rect 1975 -1355 2025 -1330
rect 2075 -1310 2125 -1300
rect 2075 -1330 2090 -1310
rect 2110 -1330 2125 -1310
rect 2075 -1355 2125 -1330
rect 2175 -1310 2225 -1300
rect 2175 -1330 2190 -1310
rect 2210 -1330 2225 -1310
rect 2175 -1355 2225 -1330
rect 2275 -1310 2325 -1300
rect 2275 -1330 2290 -1310
rect 2310 -1330 2325 -1310
rect 2665 -1320 2675 -1300
rect 2695 -1320 2720 -1300
rect 2665 -1330 2720 -1320
rect 2275 -1355 2325 -1330
rect 2375 -1355 2425 -1340
rect 2670 -1355 2720 -1330
rect 3970 -1300 4025 -1290
rect 3970 -1320 3995 -1300
rect 4015 -1320 4025 -1300
rect 3970 -1330 4025 -1320
rect 2770 -1355 2820 -1335
rect 2870 -1355 2920 -1335
rect 2970 -1355 3020 -1335
rect 3070 -1355 3120 -1335
rect 3170 -1355 3220 -1335
rect 3270 -1355 3320 -1335
rect 3370 -1355 3420 -1335
rect 3470 -1355 3520 -1335
rect 3570 -1355 3620 -1335
rect 3670 -1355 3720 -1335
rect 3770 -1355 3820 -1335
rect 3870 -1355 3920 -1335
rect 3970 -1355 4020 -1330
rect 845 -2575 895 -2555
rect 845 -2595 855 -2575
rect 875 -2595 895 -2575
rect 1075 -2580 1125 -2555
rect 1175 -2575 1225 -2555
rect 1275 -2575 1325 -2555
rect 1375 -2575 1425 -2555
rect 1475 -2575 1525 -2555
rect 1575 -2575 1625 -2555
rect 1675 -2575 1725 -2555
rect 1775 -2575 1825 -2555
rect 1875 -2575 1925 -2555
rect 1975 -2575 2025 -2555
rect 2075 -2575 2125 -2555
rect 2175 -2575 2225 -2555
rect 2275 -2575 2325 -2555
rect 845 -2605 895 -2595
rect 1070 -2590 1125 -2580
rect 1070 -2610 1080 -2590
rect 1100 -2610 1125 -2590
rect 1070 -2620 1125 -2610
rect 2375 -2580 2425 -2555
rect 2670 -2570 2720 -2555
rect 2770 -2580 2820 -2555
rect 2375 -2590 2430 -2580
rect 2375 -2610 2400 -2590
rect 2420 -2610 2430 -2590
rect 2770 -2600 2785 -2580
rect 2805 -2600 2820 -2580
rect 2770 -2610 2820 -2600
rect 2870 -2580 2920 -2555
rect 2870 -2600 2885 -2580
rect 2905 -2600 2920 -2580
rect 2870 -2610 2920 -2600
rect 2970 -2580 3020 -2555
rect 2970 -2600 2985 -2580
rect 3005 -2600 3020 -2580
rect 2970 -2610 3020 -2600
rect 3070 -2580 3120 -2555
rect 3070 -2600 3085 -2580
rect 3105 -2600 3120 -2580
rect 3070 -2610 3120 -2600
rect 3170 -2580 3220 -2555
rect 3170 -2600 3185 -2580
rect 3205 -2600 3220 -2580
rect 3170 -2610 3220 -2600
rect 3270 -2580 3320 -2555
rect 3270 -2600 3285 -2580
rect 3305 -2600 3320 -2580
rect 3270 -2610 3320 -2600
rect 3370 -2580 3420 -2555
rect 3370 -2600 3385 -2580
rect 3405 -2600 3420 -2580
rect 3370 -2610 3420 -2600
rect 3470 -2580 3520 -2555
rect 3470 -2600 3485 -2580
rect 3505 -2600 3520 -2580
rect 3470 -2610 3520 -2600
rect 3570 -2580 3620 -2555
rect 3570 -2600 3585 -2580
rect 3605 -2600 3620 -2580
rect 3570 -2610 3620 -2600
rect 3670 -2580 3720 -2555
rect 3670 -2600 3685 -2580
rect 3705 -2600 3720 -2580
rect 3670 -2610 3720 -2600
rect 3770 -2580 3820 -2555
rect 3770 -2600 3785 -2580
rect 3805 -2600 3820 -2580
rect 3770 -2610 3820 -2600
rect 3870 -2580 3920 -2555
rect 3970 -2570 4020 -2555
rect 3870 -2600 3885 -2580
rect 3905 -2600 3920 -2580
rect 3870 -2610 3920 -2600
rect 2375 -2620 2430 -2610
<< polycont >>
rect 1190 170 1210 190
rect 1290 170 1310 190
rect 1390 170 1410 190
rect 1490 170 1510 190
rect 1590 170 1610 190
rect 1690 170 1710 190
rect 1790 170 1810 190
rect 1890 170 1910 190
rect 1990 170 2010 190
rect 2090 170 2110 190
rect 2190 170 2210 190
rect 2290 170 2310 190
rect 560 55 580 75
rect 560 -45 580 -25
rect 560 -145 580 -125
rect 560 -245 580 -225
rect 560 -345 580 -325
rect 560 -445 580 -425
rect 560 -545 580 -525
rect 560 -645 580 -625
rect 560 -755 580 -735
rect 560 -845 580 -825
rect 2675 115 2695 135
rect 3995 115 4015 135
rect 1080 -1110 1100 -1090
rect 2400 -1110 2420 -1090
rect 2785 -1165 2805 -1145
rect 2885 -1165 2905 -1145
rect 2985 -1165 3005 -1145
rect 3085 -1165 3105 -1145
rect 3185 -1165 3205 -1145
rect 3285 -1165 3305 -1145
rect 3385 -1165 3405 -1145
rect 3485 -1165 3505 -1145
rect 3585 -1165 3605 -1145
rect 3685 -1165 3705 -1145
rect 3785 -1165 3805 -1145
rect 3885 -1165 3905 -1145
rect 1190 -1330 1210 -1310
rect 1290 -1330 1310 -1310
rect 1390 -1330 1410 -1310
rect 1490 -1330 1510 -1310
rect 1590 -1330 1610 -1310
rect 1690 -1330 1710 -1310
rect 1790 -1330 1810 -1310
rect 1890 -1330 1910 -1310
rect 1990 -1330 2010 -1310
rect 2090 -1330 2110 -1310
rect 2190 -1330 2210 -1310
rect 2290 -1330 2310 -1310
rect 2675 -1320 2695 -1300
rect 3995 -1320 4015 -1300
rect 855 -2595 875 -2575
rect 1080 -2610 1100 -2590
rect 2400 -2610 2420 -2590
rect 2785 -2600 2805 -2580
rect 2885 -2600 2905 -2580
rect 2985 -2600 3005 -2580
rect 3085 -2600 3105 -2580
rect 3185 -2600 3205 -2580
rect 3285 -2600 3305 -2580
rect 3385 -2600 3405 -2580
rect 3485 -2600 3505 -2580
rect 3585 -2600 3605 -2580
rect 3685 -2600 3705 -2580
rect 3785 -2600 3805 -2580
rect 3885 -2600 3905 -2580
<< locali >>
rect 920 190 2320 200
rect 610 170 900 180
rect 610 150 620 170
rect 890 150 900 170
rect 610 125 900 150
rect 610 105 620 125
rect 890 105 900 125
rect 610 95 900 105
rect 920 170 1190 190
rect 1210 170 1290 190
rect 1310 170 1390 190
rect 1410 170 1490 190
rect 1510 170 1590 190
rect 1610 170 1690 190
rect 1710 170 1790 190
rect 1810 170 1890 190
rect 1910 170 1990 190
rect 2010 170 2090 190
rect 2110 170 2190 190
rect 2210 170 2290 190
rect 2310 170 2320 190
rect 920 160 2320 170
rect 2725 160 3965 200
rect 550 75 590 85
rect 550 55 560 75
rect 580 55 590 75
rect 550 45 590 55
rect 920 35 960 160
rect 610 25 960 35
rect 610 5 620 25
rect 890 5 960 25
rect 610 -5 960 5
rect 550 -25 590 -15
rect 550 -45 560 -25
rect 580 -45 590 -25
rect 550 -125 590 -45
rect 610 -75 900 -65
rect 610 -95 620 -75
rect 890 -95 900 -75
rect 610 -105 900 -95
rect 550 -145 560 -125
rect 580 -145 590 -125
rect 550 -165 590 -145
rect 550 -175 900 -165
rect 550 -195 620 -175
rect 890 -195 900 -175
rect 550 -205 900 -195
rect 550 -225 590 -205
rect 550 -245 560 -225
rect 580 -245 590 -225
rect 550 -325 590 -245
rect 610 -275 900 -265
rect 610 -295 620 -275
rect 890 -295 900 -275
rect 610 -305 900 -295
rect 550 -345 560 -325
rect 580 -345 590 -325
rect 550 -425 590 -345
rect 920 -365 960 -5
rect 610 -375 960 -365
rect 610 -395 620 -375
rect 890 -395 960 -375
rect 610 -405 960 -395
rect 550 -445 560 -425
rect 580 -445 590 -425
rect 550 -525 590 -445
rect 610 -475 900 -465
rect 610 -495 620 -475
rect 890 -495 900 -475
rect 610 -505 900 -495
rect 550 -545 560 -525
rect 580 -545 590 -525
rect 550 -565 590 -545
rect 550 -575 900 -565
rect 550 -595 620 -575
rect 890 -595 900 -575
rect 550 -605 900 -595
rect 550 -625 590 -605
rect 550 -645 560 -625
rect 580 -645 590 -625
rect 550 -735 590 -645
rect 610 -675 900 -665
rect 610 -695 620 -675
rect 890 -695 900 -675
rect 610 -705 900 -695
rect 550 -755 560 -735
rect 580 -755 590 -735
rect 550 -765 590 -755
rect 920 -765 960 -405
rect 610 -775 960 -765
rect 610 -795 620 -775
rect 890 -795 960 -775
rect 610 -805 960 -795
rect 550 -825 590 -815
rect 550 -845 560 -825
rect 580 -845 590 -825
rect 550 -855 590 -845
rect 610 -875 900 -865
rect 610 -895 620 -875
rect 890 -895 900 -875
rect 610 -925 900 -895
rect 610 -945 620 -925
rect 890 -945 900 -925
rect 610 -955 900 -945
rect 920 -1300 960 -805
rect 980 130 1070 140
rect 980 -1040 990 130
rect 1010 -1040 1040 130
rect 1060 -1040 1070 130
rect 980 -1050 1070 -1040
rect 1130 130 1170 140
rect 1130 -1040 1140 130
rect 1160 -1040 1170 130
rect 1070 -1090 1110 -1080
rect 1070 -1110 1080 -1090
rect 1100 -1110 1110 -1090
rect 1070 -1120 1110 -1110
rect 800 -1340 960 -1300
rect 1130 -1300 1170 -1040
rect 1230 130 1270 140
rect 1230 -1040 1240 130
rect 1260 -1040 1270 130
rect 1230 -1050 1270 -1040
rect 1330 130 1370 140
rect 1330 -1040 1340 130
rect 1360 -1040 1370 130
rect 1330 -1050 1370 -1040
rect 1430 130 1470 140
rect 1430 -1040 1440 130
rect 1460 -1040 1470 130
rect 1430 -1050 1470 -1040
rect 1530 130 1570 140
rect 1530 -1040 1540 130
rect 1560 -1040 1570 130
rect 1530 -1050 1570 -1040
rect 1630 130 1670 140
rect 1630 -1040 1640 130
rect 1660 -1040 1670 130
rect 1630 -1050 1670 -1040
rect 1730 130 1770 140
rect 1730 -1040 1740 130
rect 1760 -1040 1770 130
rect 1730 -1300 1770 -1040
rect 1830 130 1870 140
rect 1830 -1040 1840 130
rect 1860 -1040 1870 130
rect 1830 -1050 1870 -1040
rect 1930 130 1970 140
rect 1930 -1040 1940 130
rect 1960 -1040 1970 130
rect 1930 -1050 1970 -1040
rect 2030 130 2070 140
rect 2030 -1040 2040 130
rect 2060 -1040 2070 130
rect 2030 -1050 2070 -1040
rect 2130 130 2170 140
rect 2130 -1040 2140 130
rect 2160 -1040 2170 130
rect 2130 -1050 2170 -1040
rect 2230 130 2270 140
rect 2230 -1040 2240 130
rect 2260 -1040 2270 130
rect 2230 -1050 2270 -1040
rect 2330 130 2370 140
rect 2330 -1040 2340 130
rect 2360 -1040 2370 130
rect 2330 -1300 2370 -1040
rect 2430 130 2515 140
rect 2430 -1040 2440 130
rect 2460 -1040 2485 130
rect 2505 -1040 2515 130
rect 2665 135 2705 145
rect 2665 115 2675 135
rect 2695 115 2705 135
rect 2665 105 2705 115
rect 2430 -1050 2515 -1040
rect 2580 65 2665 75
rect 2390 -1090 2430 -1080
rect 2390 -1110 2400 -1090
rect 2420 -1110 2430 -1090
rect 2390 -1120 2430 -1110
rect 2580 -1105 2590 65
rect 2610 -1105 2635 65
rect 2655 -1105 2665 65
rect 2580 -1115 2665 -1105
rect 2725 65 2765 160
rect 2725 -1105 2735 65
rect 2755 -1105 2765 65
rect 2725 -1135 2765 -1105
rect 2825 100 3865 140
rect 2825 65 2865 100
rect 2825 -1105 2835 65
rect 2855 -1105 2865 65
rect 2825 -1115 2865 -1105
rect 2925 65 2965 75
rect 2925 -1105 2935 65
rect 2955 -1105 2965 65
rect 2925 -1135 2965 -1105
rect 3025 65 3065 100
rect 3025 -1105 3035 65
rect 3055 -1105 3065 65
rect 3025 -1115 3065 -1105
rect 3125 65 3165 75
rect 3125 -1105 3135 65
rect 3155 -1105 3165 65
rect 3125 -1135 3165 -1105
rect 3225 65 3265 100
rect 3225 -1105 3235 65
rect 3255 -1105 3265 65
rect 3225 -1115 3265 -1105
rect 3325 65 3365 75
rect 3325 -1105 3335 65
rect 3355 -1105 3365 65
rect 3325 -1115 3365 -1105
rect 3425 65 3465 100
rect 3425 -1105 3435 65
rect 3455 -1105 3465 65
rect 3425 -1115 3465 -1105
rect 3525 65 3565 75
rect 3525 -1105 3535 65
rect 3555 -1105 3565 65
rect 3525 -1135 3565 -1105
rect 3625 65 3665 100
rect 3625 -1105 3635 65
rect 3655 -1105 3665 65
rect 3625 -1115 3665 -1105
rect 3725 65 3765 75
rect 3725 -1105 3735 65
rect 3755 -1105 3765 65
rect 3725 -1135 3765 -1105
rect 3825 65 3865 100
rect 3825 -1105 3835 65
rect 3855 -1105 3865 65
rect 3825 -1115 3865 -1105
rect 3925 65 3965 160
rect 3985 135 4025 145
rect 3985 115 3995 135
rect 4015 115 4025 135
rect 3985 105 4025 115
rect 3925 -1105 3935 65
rect 3955 -1105 3965 65
rect 3925 -1135 3965 -1105
rect 4025 65 4115 75
rect 4025 -1105 4035 65
rect 4055 -1105 4085 65
rect 4105 -1105 4115 65
rect 4025 -1115 4115 -1105
rect 2725 -1145 2815 -1135
rect 2725 -1165 2785 -1145
rect 2805 -1165 2815 -1145
rect 2725 -1175 2815 -1165
rect 2875 -1145 3815 -1135
rect 2875 -1165 2885 -1145
rect 2905 -1165 2985 -1145
rect 3005 -1165 3085 -1145
rect 3105 -1165 3185 -1145
rect 3205 -1165 3285 -1145
rect 3305 -1165 3385 -1145
rect 3405 -1165 3485 -1145
rect 3505 -1165 3585 -1145
rect 3605 -1165 3685 -1145
rect 3705 -1165 3785 -1145
rect 3805 -1165 3815 -1145
rect 2875 -1175 3815 -1165
rect 3875 -1145 3965 -1135
rect 3875 -1165 3885 -1145
rect 3905 -1165 3965 -1145
rect 3875 -1175 3965 -1165
rect 1130 -1310 1220 -1300
rect 1130 -1330 1190 -1310
rect 1210 -1330 1220 -1310
rect 1130 -1340 1220 -1330
rect 1280 -1310 2220 -1300
rect 1280 -1330 1290 -1310
rect 1310 -1330 1390 -1310
rect 1410 -1330 1490 -1310
rect 1510 -1330 1590 -1310
rect 1610 -1330 1690 -1310
rect 1710 -1330 1790 -1310
rect 1810 -1330 1890 -1310
rect 1910 -1330 1990 -1310
rect 2010 -1330 2090 -1310
rect 2110 -1330 2190 -1310
rect 2210 -1330 2220 -1310
rect 1280 -1340 2220 -1330
rect 2280 -1310 2370 -1300
rect 2280 -1330 2290 -1310
rect 2310 -1330 2370 -1310
rect 2665 -1300 2705 -1290
rect 2665 -1320 2675 -1300
rect 2695 -1320 2705 -1300
rect 2665 -1330 2705 -1320
rect 2280 -1340 2370 -1330
rect 800 -1370 840 -1340
rect 800 -2535 810 -1370
rect 830 -2535 840 -1370
rect 800 -2565 840 -2535
rect 900 -1370 940 -1360
rect 900 -2535 910 -1370
rect 930 -2535 940 -1370
rect 900 -2550 940 -2535
rect 980 -1370 1070 -1360
rect 980 -2540 990 -1370
rect 1010 -2540 1040 -1370
rect 1060 -2540 1070 -1370
rect 980 -2550 1070 -2540
rect 1130 -1370 1170 -1340
rect 1130 -2540 1140 -1370
rect 1160 -2540 1170 -1370
rect 800 -2575 885 -2565
rect 800 -2595 855 -2575
rect 875 -2595 885 -2575
rect 800 -2605 885 -2595
rect 1070 -2590 1110 -2580
rect 1070 -2610 1080 -2590
rect 1100 -2610 1110 -2590
rect 1070 -2620 1110 -2610
rect 1130 -2635 1170 -2540
rect 1230 -1370 1270 -1360
rect 1230 -2540 1240 -1370
rect 1260 -2540 1270 -1370
rect 1230 -2575 1270 -2540
rect 1330 -1370 1370 -1340
rect 1330 -2540 1340 -1370
rect 1360 -2540 1370 -1370
rect 1330 -2550 1370 -2540
rect 1430 -1370 1470 -1360
rect 1430 -2540 1440 -1370
rect 1460 -2540 1470 -1370
rect 1430 -2575 1470 -2540
rect 1530 -1370 1570 -1340
rect 1530 -2540 1540 -1370
rect 1560 -2540 1570 -1370
rect 1530 -2550 1570 -2540
rect 1630 -1370 1670 -1360
rect 1630 -2540 1640 -1370
rect 1660 -2540 1670 -1370
rect 1630 -2575 1670 -2540
rect 1730 -1370 1770 -1360
rect 1730 -2540 1740 -1370
rect 1760 -2540 1770 -1370
rect 1730 -2550 1770 -2540
rect 1830 -1370 1870 -1360
rect 1830 -2540 1840 -1370
rect 1860 -2540 1870 -1370
rect 1830 -2575 1870 -2540
rect 1930 -1370 1970 -1340
rect 1930 -2540 1940 -1370
rect 1960 -2540 1970 -1370
rect 1930 -2550 1970 -2540
rect 2030 -1370 2070 -1360
rect 2030 -2540 2040 -1370
rect 2060 -2540 2070 -1370
rect 2030 -2575 2070 -2540
rect 2130 -1370 2170 -1340
rect 2130 -2540 2140 -1370
rect 2160 -2540 2170 -1370
rect 2130 -2550 2170 -2540
rect 2230 -1370 2270 -1360
rect 2230 -2540 2240 -1370
rect 2260 -2540 2270 -1370
rect 2230 -2575 2270 -2540
rect 1230 -2615 2270 -2575
rect 2330 -1370 2370 -1340
rect 2330 -2540 2340 -1370
rect 2360 -2540 2370 -1370
rect 2330 -2635 2370 -2540
rect 2430 -1370 2515 -1360
rect 2430 -2540 2440 -1370
rect 2460 -2540 2485 -1370
rect 2505 -2540 2515 -1370
rect 2430 -2550 2515 -2540
rect 2580 -1370 2665 -1360
rect 2580 -2540 2590 -1370
rect 2610 -2540 2635 -1370
rect 2655 -2540 2665 -1370
rect 2580 -2550 2665 -2540
rect 2725 -1370 2765 -1175
rect 2725 -2540 2735 -1370
rect 2755 -2540 2765 -1370
rect 2725 -2550 2765 -2540
rect 2825 -1370 2865 -1360
rect 2825 -2540 2835 -1370
rect 2855 -2540 2865 -1370
rect 2825 -2550 2865 -2540
rect 2925 -1370 2965 -1360
rect 2925 -2540 2935 -1370
rect 2955 -2540 2965 -1370
rect 2925 -2550 2965 -2540
rect 3025 -1370 3065 -1360
rect 3025 -2540 3035 -1370
rect 3055 -2540 3065 -1370
rect 3025 -2550 3065 -2540
rect 3125 -1370 3165 -1360
rect 3125 -2540 3135 -1370
rect 3155 -2540 3165 -1370
rect 3125 -2550 3165 -2540
rect 3225 -1370 3265 -1360
rect 3225 -2540 3235 -1370
rect 3255 -2540 3265 -1370
rect 3225 -2550 3265 -2540
rect 3325 -1370 3365 -1175
rect 3325 -2540 3335 -1370
rect 3355 -2540 3365 -1370
rect 3325 -2550 3365 -2540
rect 3425 -1370 3465 -1360
rect 3425 -2540 3435 -1370
rect 3455 -2540 3465 -1370
rect 3425 -2550 3465 -2540
rect 3525 -1370 3565 -1360
rect 3525 -2540 3535 -1370
rect 3555 -2540 3565 -1370
rect 3525 -2550 3565 -2540
rect 3625 -1370 3665 -1360
rect 3625 -2540 3635 -1370
rect 3655 -2540 3665 -1370
rect 3625 -2550 3665 -2540
rect 3725 -1370 3765 -1360
rect 3725 -2540 3735 -1370
rect 3755 -2540 3765 -1370
rect 3725 -2550 3765 -2540
rect 3825 -1370 3865 -1360
rect 3825 -2540 3835 -1370
rect 3855 -2540 3865 -1370
rect 3825 -2550 3865 -2540
rect 3925 -1370 3965 -1175
rect 3985 -1300 4025 -1290
rect 3985 -1320 3995 -1300
rect 4015 -1320 4025 -1300
rect 3985 -1330 4025 -1320
rect 3925 -2540 3935 -1370
rect 3955 -2540 3965 -1370
rect 3925 -2550 3965 -2540
rect 4025 -1370 4115 -1360
rect 4025 -2540 4035 -1370
rect 4055 -2540 4085 -1370
rect 4105 -2540 4115 -1370
rect 4025 -2550 4115 -2540
rect 2775 -2580 3915 -2570
rect 2390 -2590 2430 -2580
rect 2390 -2610 2400 -2590
rect 2420 -2610 2430 -2590
rect 2775 -2600 2785 -2580
rect 2805 -2600 2885 -2580
rect 2905 -2600 2985 -2580
rect 3005 -2600 3085 -2580
rect 3105 -2600 3185 -2580
rect 3205 -2600 3285 -2580
rect 3305 -2600 3385 -2580
rect 3405 -2600 3485 -2580
rect 3505 -2600 3585 -2580
rect 3605 -2600 3685 -2580
rect 3705 -2600 3785 -2580
rect 3805 -2600 3885 -2580
rect 3905 -2600 3915 -2580
rect 2775 -2610 3915 -2600
rect 2390 -2620 2430 -2610
rect 1130 -2675 2370 -2635
<< viali >>
rect 620 150 890 170
rect 620 105 890 125
rect 560 55 580 75
rect 620 -95 890 -75
rect 620 -295 890 -275
rect 620 -495 890 -475
rect 620 -695 890 -675
rect 560 -845 580 -825
rect 620 -895 890 -875
rect 620 -945 890 -925
rect 990 -1040 1010 130
rect 1040 -1040 1060 130
rect 1240 -1040 1260 130
rect 2240 -1040 2260 130
rect 2440 -1040 2460 130
rect 2485 -1040 2505 130
rect 2590 -1105 2610 65
rect 2635 -1105 2655 65
rect 3335 -1105 3355 65
rect 4035 -1105 4055 65
rect 4085 -1105 4105 65
rect 910 -2535 930 -1370
rect 990 -2540 1010 -1370
rect 1040 -2540 1060 -1370
rect 1740 -2540 1760 -1370
rect 2440 -2540 2460 -1370
rect 2485 -2540 2505 -1370
rect 2590 -2540 2610 -1370
rect 2635 -2540 2655 -1370
rect 2835 -2540 2855 -1370
rect 3835 -2540 3855 -1370
rect 4035 -2540 4055 -1370
rect 4085 -2540 4105 -1370
<< metal1 >>
rect 610 170 900 180
rect 610 150 620 170
rect 890 150 900 170
rect 610 140 900 150
rect 610 130 2515 140
rect 610 125 990 130
rect 610 105 620 125
rect 890 105 990 125
rect 610 85 990 105
rect 550 75 990 85
rect 550 55 560 75
rect 580 55 990 75
rect 550 45 990 55
rect 610 -75 990 45
rect 610 -95 620 -75
rect 890 -95 990 -75
rect 610 -275 990 -95
rect 610 -295 620 -275
rect 890 -295 990 -275
rect 610 -475 990 -295
rect 610 -495 620 -475
rect 890 -495 990 -475
rect 610 -675 990 -495
rect 610 -695 620 -675
rect 890 -695 990 -675
rect 610 -705 990 -695
rect 625 -765 990 -705
rect 610 -815 990 -765
rect 550 -825 990 -815
rect 550 -845 560 -825
rect 580 -845 990 -825
rect 550 -855 990 -845
rect 610 -875 990 -855
rect 610 -895 620 -875
rect 890 -895 990 -875
rect 610 -925 990 -895
rect 610 -945 620 -925
rect 890 -945 990 -925
rect 610 -955 990 -945
rect 980 -1040 990 -955
rect 1010 -1040 1040 130
rect 1060 -1040 1240 130
rect 1260 -1040 2240 130
rect 2260 -1040 2440 130
rect 2460 -1040 2485 130
rect 2505 75 2515 130
rect 2665 105 2720 145
rect 2670 75 2720 105
rect 3970 105 4025 145
rect 3970 75 4020 105
rect 2505 65 4115 75
rect 2505 -1040 2590 65
rect 980 -1050 2590 -1040
rect 1075 -1080 1125 -1050
rect 1070 -1120 1125 -1080
rect 2375 -1080 2425 -1050
rect 2375 -1120 2430 -1080
rect 2580 -1105 2590 -1050
rect 2610 -1105 2635 65
rect 2655 -1105 3335 65
rect 3355 -1105 4035 65
rect 4055 -1105 4085 65
rect 4105 -1105 4115 65
rect 2580 -1115 4115 -1105
rect 2665 -1330 2720 -1290
rect 2670 -1360 2720 -1330
rect 3970 -1330 4025 -1290
rect 3970 -1360 4020 -1330
rect 900 -1370 4115 -1360
rect 900 -2535 910 -1370
rect 930 -2535 990 -1370
rect 900 -2540 990 -2535
rect 1010 -2540 1040 -1370
rect 1060 -2540 1740 -1370
rect 1760 -2540 2440 -1370
rect 2460 -2540 2485 -1370
rect 2505 -2540 2590 -1370
rect 2610 -2540 2635 -1370
rect 2655 -2540 2835 -1370
rect 2855 -2540 3835 -1370
rect 3855 -2540 4035 -1370
rect 4055 -2540 4085 -1370
rect 4105 -2540 4115 -1370
rect 900 -2545 4115 -2540
rect 980 -2550 4115 -2545
rect 1075 -2580 1125 -2550
rect 1070 -2620 1125 -2580
rect 2375 -2580 2425 -2550
rect 2375 -2620 2430 -2580
<< labels >>
rlabel metal1 610 160 610 160 7 VP
port 1 w
rlabel metal1 920 -1360 920 -1360 1 VN
port 2 n
rlabel locali 800 -2585 800 -2585 7 VBN
port 4 w
rlabel locali 550 -745 550 -745 7 VBP
port 3 w
rlabel locali 1130 -2655 1130 -2655 7 VCN
port 5 w
rlabel locali 2795 -2610 2795 -2610 5 VCP
port 6 s
<< end >>
