magic
tech sky130A
timestamp 1695600092
<< end >>
