magic
tech sky130A
timestamp 1695849814
<< nwell >>
rect -115 125 90 265
<< nmos >>
rect 5 -95 20 5
<< pmos >>
rect 5 145 20 245
<< ndiff >>
rect -45 -10 5 5
rect -45 -80 -30 -10
rect -10 -80 5 -10
rect -45 -95 5 -80
rect 20 -10 70 5
rect 20 -80 35 -10
rect 55 -80 70 -10
rect 20 -95 70 -80
<< pdiff >>
rect -45 230 5 245
rect -45 160 -30 230
rect -10 160 5 230
rect -45 145 5 160
rect 20 230 70 245
rect 20 160 35 230
rect 55 160 70 230
rect 20 145 70 160
<< ndiffc >>
rect -30 -80 -10 -10
rect 35 -80 55 -10
<< pdiffc >>
rect -30 160 -10 230
rect 35 160 55 230
<< psubdiff >>
rect -95 -10 -45 5
rect -95 -80 -80 -10
rect -60 -80 -45 -10
rect -95 -95 -45 -80
<< nsubdiff >>
rect -95 230 -45 245
rect -95 160 -80 230
rect -60 160 -45 230
rect -95 145 -45 160
<< psubdiffcont >>
rect -80 -80 -60 -10
<< nsubdiffcont >>
rect -80 160 -60 230
<< poly >>
rect -20 290 20 300
rect -20 270 -10 290
rect 10 270 20 290
rect -20 260 20 270
rect 5 245 20 260
rect 5 5 20 145
rect 5 -110 20 -95
<< polycont >>
rect -10 270 10 290
<< locali >>
rect -20 290 20 300
rect -20 280 -10 290
rect -115 270 -10 280
rect 10 270 20 290
rect -115 260 20 270
rect -90 230 0 240
rect -90 160 -80 230
rect -60 160 -30 230
rect -10 160 0 230
rect -90 150 0 160
rect 25 230 65 240
rect 25 160 35 230
rect 55 220 65 230
rect 55 200 90 220
rect 55 160 65 200
rect 25 150 65 160
rect 45 0 65 150
rect -90 -10 0 0
rect -90 -80 -80 -10
rect -60 -80 -30 -10
rect -10 -80 0 -10
rect -90 -90 0 -80
rect 25 -10 65 0
rect 25 -80 35 -10
rect 55 -80 65 -10
rect 25 -90 65 -80
<< viali >>
rect -80 160 -60 230
rect -30 160 -10 230
rect -80 -80 -60 -10
rect -30 -80 -10 -10
<< metal1 >>
rect -95 230 70 245
rect -95 160 -80 230
rect -60 160 -30 230
rect -10 160 70 230
rect -95 145 70 160
rect -95 -10 70 5
rect -95 -80 -80 -10
rect -60 -80 -30 -10
rect -10 -80 70 -10
rect -95 -95 70 -80
<< labels >>
rlabel locali -115 270 -115 270 7 A
port 1 w
rlabel locali 90 210 90 210 3 Y
port 2 e
rlabel metal1 -95 -45 -95 -45 7 VN
port 4 w
rlabel metal1 -95 195 -95 195 7 VP
port 3 w
<< end >>
