magic
tech sky130A
timestamp 1697389794
<< nwell >>
rect -7020 1705 -6970 2895
<< poly >>
rect -6780 145 -6740 155
rect -6655 145 -6615 155
rect -6780 125 -6770 145
rect -6750 130 -6645 145
rect -6750 125 -6740 130
rect -6780 115 -6740 125
rect -6655 125 -6645 130
rect -6625 125 -6615 145
rect -6655 115 -6615 125
<< polycont >>
rect -6770 125 -6750 145
rect -6645 125 -6625 145
<< locali >>
rect -8830 2890 -8230 2930
rect -8830 155 -8790 2890
rect -8270 2680 -8230 2890
rect -7660 2910 -4755 2950
rect -7660 2680 -7620 2910
rect -4795 2890 -4755 2910
rect -8275 2640 -8230 2680
rect -7675 2640 -7620 2680
rect -7025 1930 -6970 1975
rect -7950 225 -7910 465
rect -7950 185 -6720 225
rect -8830 145 -6740 155
rect -8830 125 -6770 145
rect -6750 125 -6740 145
rect -8830 115 -6740 125
rect -6655 150 -6465 155
rect -6390 150 -6380 155
rect -6655 145 -6380 150
rect -6655 125 -6645 145
rect -6625 125 -6380 145
rect -6655 115 -6380 125
<< metal1 >>
rect -7100 1730 -6910 2830
rect -7200 390 -6620 1460
use bias_generator  bias_generator_0
timestamp 1697389219
transform 1 0 -7520 0 1 2690
box 550 -2635 4140 205
use folded_cascode_differential_amplifier  folded_cascode_differential_amplifier_0 ~/Documents/VLSI/mp3/layouts
timestamp 1697388805
transform 0 1 -7190 -1 0 2785
box -110 -1580 2410 170
<< end >>
