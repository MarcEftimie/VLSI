magic
tech sky130A
timestamp 1697321830
<< nwell >>
rect -110 -230 1080 170
rect -110 -480 1085 -230
rect -110 -880 1240 -480
<< nmos >>
rect 1350 -305 1400 -5
rect 1450 -305 1500 -5
rect 1550 -305 1600 -5
rect 1650 -305 1700 -5
rect 1750 -305 1800 -5
rect 1850 -305 1900 -5
rect 1950 -305 2000 -5
rect 2050 -305 2100 -5
rect 2150 -305 2200 -5
rect 2250 -305 2300 -5
rect 1605 -660 2205 -610
rect 1605 -760 2205 -710
rect 10 -1455 60 -1155
rect 110 -1455 160 -1155
rect 210 -1455 260 -1155
rect 390 -1455 440 -1155
rect 490 -1455 540 -1155
rect 590 -1455 640 -1155
rect 690 -1455 740 -1155
rect 870 -1455 920 -1155
rect 970 -1455 1020 -1155
rect 1070 -1455 1120 -1155
rect 1350 -1375 1400 -1075
rect 1450 -1375 1500 -1075
rect 1550 -1375 1600 -1075
rect 1655 -1375 1705 -1075
rect 1755 -1375 1805 -1075
rect 1855 -1375 1905 -1075
rect 1955 -1375 2005 -1075
rect 2060 -1375 2110 -1075
rect 2160 -1375 2210 -1075
rect 2260 -1375 2310 -1075
<< pmos >>
rect 10 -205 60 95
rect 110 -205 160 95
rect 210 -205 260 95
rect 310 -205 360 95
rect 410 -205 460 95
rect 510 -205 560 95
rect 610 -205 660 95
rect 710 -205 760 95
rect 810 -205 860 95
rect 910 -205 960 95
rect 10 -855 60 -555
rect 110 -855 160 -555
rect 210 -855 260 -555
rect 390 -855 440 -555
rect 490 -855 540 -555
rect 590 -855 640 -555
rect 690 -855 740 -555
rect 870 -855 920 -555
rect 970 -855 1020 -555
rect 1070 -855 1120 -555
<< ndiff >>
rect 1300 -20 1350 -5
rect 1300 -290 1315 -20
rect 1335 -290 1350 -20
rect 1300 -305 1350 -290
rect 1400 -20 1450 -5
rect 1400 -290 1415 -20
rect 1435 -290 1450 -20
rect 1400 -305 1450 -290
rect 1500 -20 1550 -5
rect 1500 -290 1515 -20
rect 1535 -290 1550 -20
rect 1500 -305 1550 -290
rect 1600 -20 1650 -5
rect 1600 -290 1615 -20
rect 1635 -290 1650 -20
rect 1600 -305 1650 -290
rect 1700 -20 1750 -5
rect 1700 -290 1715 -20
rect 1735 -290 1750 -20
rect 1700 -305 1750 -290
rect 1800 -20 1850 -5
rect 1800 -290 1815 -20
rect 1835 -290 1850 -20
rect 1800 -305 1850 -290
rect 1900 -20 1950 -5
rect 1900 -290 1915 -20
rect 1935 -290 1950 -20
rect 1900 -305 1950 -290
rect 2000 -20 2050 -5
rect 2000 -290 2015 -20
rect 2035 -290 2050 -20
rect 2000 -305 2050 -290
rect 2100 -20 2150 -5
rect 2100 -290 2115 -20
rect 2135 -290 2150 -20
rect 2100 -305 2150 -290
rect 2200 -20 2250 -5
rect 2200 -290 2215 -20
rect 2235 -290 2250 -20
rect 2200 -305 2250 -290
rect 2300 -20 2350 -5
rect 2300 -290 2315 -20
rect 2335 -290 2350 -20
rect 2300 -305 2350 -290
rect 1605 -575 2205 -560
rect 1605 -595 1620 -575
rect 2190 -595 2205 -575
rect 1605 -610 2205 -595
rect 1605 -675 2205 -660
rect 1605 -695 1620 -675
rect 2190 -695 2205 -675
rect 1605 -710 2205 -695
rect 1605 -775 2205 -760
rect 1605 -795 1620 -775
rect 2190 -795 2205 -775
rect 1605 -810 2205 -795
rect -40 -1170 10 -1155
rect -40 -1440 -25 -1170
rect -5 -1440 10 -1170
rect -40 -1455 10 -1440
rect 60 -1170 110 -1155
rect 60 -1440 75 -1170
rect 95 -1440 110 -1170
rect 60 -1455 110 -1440
rect 160 -1170 210 -1155
rect 160 -1440 175 -1170
rect 195 -1440 210 -1170
rect 160 -1455 210 -1440
rect 260 -1170 310 -1155
rect 260 -1440 275 -1170
rect 295 -1440 310 -1170
rect 260 -1455 310 -1440
rect 340 -1170 390 -1155
rect 340 -1440 355 -1170
rect 375 -1440 390 -1170
rect 340 -1455 390 -1440
rect 440 -1170 490 -1155
rect 440 -1440 455 -1170
rect 475 -1440 490 -1170
rect 440 -1455 490 -1440
rect 540 -1170 590 -1155
rect 540 -1440 555 -1170
rect 575 -1440 590 -1170
rect 540 -1455 590 -1440
rect 640 -1170 690 -1155
rect 640 -1440 655 -1170
rect 675 -1440 690 -1170
rect 640 -1455 690 -1440
rect 740 -1170 790 -1155
rect 740 -1440 755 -1170
rect 775 -1440 790 -1170
rect 740 -1455 790 -1440
rect 820 -1170 870 -1155
rect 820 -1440 835 -1170
rect 855 -1440 870 -1170
rect 820 -1455 870 -1440
rect 920 -1170 970 -1155
rect 920 -1440 935 -1170
rect 955 -1440 970 -1170
rect 920 -1455 970 -1440
rect 1020 -1170 1070 -1155
rect 1020 -1440 1035 -1170
rect 1055 -1440 1070 -1170
rect 1020 -1455 1070 -1440
rect 1120 -1170 1170 -1155
rect 1120 -1440 1135 -1170
rect 1155 -1440 1170 -1170
rect 1120 -1455 1170 -1440
rect 1300 -1090 1350 -1075
rect 1300 -1360 1315 -1090
rect 1335 -1360 1350 -1090
rect 1300 -1375 1350 -1360
rect 1400 -1090 1450 -1075
rect 1400 -1360 1415 -1090
rect 1435 -1360 1450 -1090
rect 1400 -1375 1450 -1360
rect 1500 -1090 1550 -1075
rect 1500 -1360 1515 -1090
rect 1535 -1360 1550 -1090
rect 1500 -1375 1550 -1360
rect 1600 -1090 1655 -1075
rect 1600 -1360 1620 -1090
rect 1640 -1360 1655 -1090
rect 1600 -1375 1655 -1360
rect 1705 -1090 1755 -1075
rect 1705 -1360 1720 -1090
rect 1740 -1360 1755 -1090
rect 1705 -1375 1755 -1360
rect 1805 -1090 1855 -1075
rect 1805 -1360 1820 -1090
rect 1840 -1360 1855 -1090
rect 1805 -1375 1855 -1360
rect 1905 -1090 1955 -1075
rect 1905 -1360 1920 -1090
rect 1940 -1360 1955 -1090
rect 1905 -1375 1955 -1360
rect 2005 -1090 2060 -1075
rect 2005 -1360 2025 -1090
rect 2045 -1360 2060 -1090
rect 2005 -1375 2060 -1360
rect 2110 -1090 2160 -1075
rect 2110 -1360 2125 -1090
rect 2145 -1360 2160 -1090
rect 2110 -1375 2160 -1360
rect 2210 -1090 2260 -1075
rect 2210 -1360 2225 -1090
rect 2245 -1360 2260 -1090
rect 2210 -1375 2260 -1360
rect 2310 -1090 2360 -1075
rect 2310 -1360 2325 -1090
rect 2345 -1360 2360 -1090
rect 2310 -1375 2360 -1360
<< pdiff >>
rect -40 80 10 95
rect -40 -190 -25 80
rect -5 -190 10 80
rect -40 -205 10 -190
rect 60 80 110 95
rect 60 -190 75 80
rect 95 -190 110 80
rect 60 -205 110 -190
rect 160 80 210 95
rect 160 -190 175 80
rect 195 -190 210 80
rect 160 -205 210 -190
rect 260 80 310 95
rect 260 -190 275 80
rect 295 -190 310 80
rect 260 -205 310 -190
rect 360 80 410 95
rect 360 -190 375 80
rect 395 -190 410 80
rect 360 -205 410 -190
rect 460 80 510 95
rect 460 -190 475 80
rect 495 -190 510 80
rect 460 -205 510 -190
rect 560 80 610 95
rect 560 -190 575 80
rect 595 -190 610 80
rect 560 -205 610 -190
rect 660 80 710 95
rect 660 -190 675 80
rect 695 -190 710 80
rect 660 -205 710 -190
rect 760 80 810 95
rect 760 -190 775 80
rect 795 -190 810 80
rect 760 -205 810 -190
rect 860 80 910 95
rect 860 -190 875 80
rect 895 -190 910 80
rect 860 -205 910 -190
rect 960 80 1010 95
rect 960 -190 975 80
rect 995 -190 1010 80
rect 960 -205 1010 -190
rect -40 -570 10 -555
rect -40 -840 -25 -570
rect -5 -840 10 -570
rect -40 -855 10 -840
rect 60 -570 110 -555
rect 60 -840 75 -570
rect 95 -840 110 -570
rect 60 -855 110 -840
rect 160 -570 210 -555
rect 160 -840 175 -570
rect 195 -840 210 -570
rect 160 -855 210 -840
rect 260 -570 310 -555
rect 260 -840 275 -570
rect 295 -840 310 -570
rect 260 -855 310 -840
rect 340 -570 390 -555
rect 340 -840 355 -570
rect 375 -840 390 -570
rect 340 -855 390 -840
rect 440 -570 490 -555
rect 440 -840 455 -570
rect 475 -840 490 -570
rect 440 -855 490 -840
rect 540 -570 590 -555
rect 540 -840 555 -570
rect 575 -840 590 -570
rect 540 -855 590 -840
rect 640 -570 690 -555
rect 640 -840 655 -570
rect 675 -840 690 -570
rect 640 -855 690 -840
rect 740 -570 790 -555
rect 740 -840 755 -570
rect 775 -840 790 -570
rect 740 -855 790 -840
rect 820 -570 870 -555
rect 820 -840 835 -570
rect 855 -840 870 -570
rect 820 -855 870 -840
rect 920 -570 970 -555
rect 920 -840 935 -570
rect 955 -840 970 -570
rect 920 -855 970 -840
rect 1020 -570 1070 -555
rect 1020 -840 1035 -570
rect 1055 -840 1070 -570
rect 1020 -855 1070 -840
rect 1120 -570 1170 -555
rect 1120 -840 1135 -570
rect 1155 -840 1170 -570
rect 1120 -855 1170 -840
<< ndiffc >>
rect 1315 -290 1335 -20
rect 1415 -290 1435 -20
rect 1515 -290 1535 -20
rect 1615 -290 1635 -20
rect 1715 -290 1735 -20
rect 1815 -290 1835 -20
rect 1915 -290 1935 -20
rect 2015 -290 2035 -20
rect 2115 -290 2135 -20
rect 2215 -290 2235 -20
rect 2315 -290 2335 -20
rect 1620 -595 2190 -575
rect 1620 -695 2190 -675
rect 1620 -795 2190 -775
rect -25 -1440 -5 -1170
rect 75 -1440 95 -1170
rect 175 -1440 195 -1170
rect 275 -1440 295 -1170
rect 355 -1440 375 -1170
rect 455 -1440 475 -1170
rect 555 -1440 575 -1170
rect 655 -1440 675 -1170
rect 755 -1440 775 -1170
rect 835 -1440 855 -1170
rect 935 -1440 955 -1170
rect 1035 -1440 1055 -1170
rect 1135 -1440 1155 -1170
rect 1315 -1360 1335 -1090
rect 1415 -1360 1435 -1090
rect 1515 -1360 1535 -1090
rect 1620 -1360 1640 -1090
rect 1720 -1360 1740 -1090
rect 1820 -1360 1840 -1090
rect 1920 -1360 1940 -1090
rect 2025 -1360 2045 -1090
rect 2125 -1360 2145 -1090
rect 2225 -1360 2245 -1090
rect 2325 -1360 2345 -1090
<< pdiffc >>
rect -25 -190 -5 80
rect 75 -190 95 80
rect 175 -190 195 80
rect 275 -190 295 80
rect 375 -190 395 80
rect 475 -190 495 80
rect 575 -190 595 80
rect 675 -190 695 80
rect 775 -190 795 80
rect 875 -190 895 80
rect 975 -190 995 80
rect -25 -840 -5 -570
rect 75 -840 95 -570
rect 175 -840 195 -570
rect 275 -840 295 -570
rect 355 -840 375 -570
rect 455 -840 475 -570
rect 555 -840 575 -570
rect 655 -840 675 -570
rect 755 -840 775 -570
rect 835 -840 855 -570
rect 935 -840 955 -570
rect 1035 -840 1055 -570
rect 1135 -840 1155 -570
<< psubdiff >>
rect 1250 -20 1300 -5
rect 1250 -290 1265 -20
rect 1285 -290 1300 -20
rect 1250 -305 1300 -290
rect 2350 -305 2400 -5
rect -90 -1170 -40 -1155
rect -90 -1365 -75 -1170
rect -55 -1365 -40 -1170
rect -90 -1455 -40 -1365
rect 1170 -1455 1220 -1155
rect 1250 -1375 1300 -1075
rect 2360 -1375 2410 -1075
<< nsubdiff >>
rect -90 80 -40 95
rect -90 -190 -75 80
rect -55 -190 -40 80
rect -90 -205 -40 -190
rect 1010 80 1060 95
rect 1010 -190 1025 80
rect 1045 -190 1060 80
rect 1010 -205 1060 -190
rect -90 -570 -40 -555
rect -90 -840 -75 -570
rect -55 -840 -40 -570
rect -90 -855 -40 -840
rect 1170 -570 1220 -555
rect 1170 -840 1185 -570
rect 1205 -840 1220 -570
rect 1170 -855 1220 -840
<< psubdiffcont >>
rect 1265 -290 1285 -20
rect -75 -1365 -55 -1170
<< nsubdiffcont >>
rect -75 -190 -55 80
rect 1025 -190 1045 80
rect -75 -840 -55 -570
rect 1185 -840 1205 -570
<< poly >>
rect 110 155 160 170
rect 10 140 60 155
rect 10 120 25 140
rect 45 120 60 140
rect 10 95 60 120
rect 110 135 125 155
rect 145 135 160 155
rect 110 95 160 135
rect 210 155 260 170
rect 210 135 225 155
rect 245 135 260 155
rect 210 95 260 135
rect 310 155 360 170
rect 310 135 325 155
rect 345 135 360 155
rect 310 95 360 135
rect 410 155 460 170
rect 410 135 425 155
rect 445 135 460 155
rect 410 95 460 135
rect 510 155 560 170
rect 510 135 525 155
rect 545 135 560 155
rect 510 95 560 135
rect 610 155 660 170
rect 610 135 625 155
rect 645 135 660 155
rect 610 95 660 135
rect 710 155 760 170
rect 710 135 725 155
rect 745 135 760 155
rect 710 95 760 135
rect 810 155 860 170
rect 810 135 825 155
rect 845 135 860 155
rect 810 95 860 135
rect 910 140 960 155
rect 910 120 925 140
rect 945 120 960 140
rect 910 95 960 120
rect 1450 45 2200 60
rect 1350 -5 1400 20
rect 1450 -5 1500 45
rect 1550 -5 1600 20
rect 1650 -5 1700 20
rect 1750 -5 1800 45
rect 1850 -5 1900 45
rect 1950 -5 2000 20
rect 2050 -5 2100 20
rect 2150 -5 2200 45
rect 2250 -5 2300 20
rect 10 -230 60 -205
rect 110 -230 160 -205
rect 210 -230 260 -205
rect 310 -230 360 -205
rect 410 -230 460 -205
rect 510 -230 560 -205
rect 610 -230 660 -205
rect 710 -230 760 -205
rect 810 -230 860 -205
rect 910 -230 960 -205
rect 405 -265 965 -255
rect 405 -285 415 -265
rect 435 -270 675 -265
rect 435 -285 445 -270
rect 405 -295 445 -285
rect 665 -285 675 -270
rect 695 -270 935 -265
rect 695 -285 705 -270
rect 665 -295 705 -285
rect 925 -285 935 -270
rect 955 -285 965 -265
rect 925 -295 965 -285
rect 1350 -325 1400 -305
rect 1450 -315 1500 -305
rect 1350 -345 1365 -325
rect 1385 -345 1400 -325
rect 1350 -360 1400 -345
rect 1445 -325 1500 -315
rect 1445 -345 1455 -325
rect 1475 -345 1500 -325
rect 1445 -355 1500 -345
rect 1550 -355 1600 -305
rect 1650 -355 1700 -305
rect 1750 -330 1800 -305
rect 1850 -330 1900 -305
rect 1950 -355 2000 -305
rect 2050 -355 2100 -305
rect 2150 -320 2200 -305
rect 1550 -370 2100 -355
rect 2250 -325 2300 -305
rect 2250 -345 2265 -325
rect 2285 -345 2300 -325
rect 2250 -360 2300 -345
rect 2080 -385 2100 -370
rect 2080 -395 2120 -385
rect 485 -405 525 -395
rect 485 -425 495 -405
rect 515 -420 525 -405
rect 605 -405 645 -395
rect 605 -420 615 -405
rect 515 -425 615 -420
rect 635 -425 645 -405
rect 485 -435 645 -425
rect 1445 -405 1485 -395
rect 1445 -425 1455 -405
rect 1475 -420 1485 -405
rect 1605 -405 1645 -395
rect 1605 -420 1615 -405
rect 1475 -425 1615 -420
rect 1635 -420 1645 -405
rect 2005 -405 2045 -395
rect 2005 -420 2015 -405
rect 1635 -425 2015 -420
rect 2035 -425 2045 -405
rect 2080 -415 2090 -395
rect 2110 -415 2120 -395
rect 2080 -425 2120 -415
rect 1445 -435 2045 -425
rect 100 -495 1020 -480
rect 10 -510 60 -495
rect 10 -530 25 -510
rect 45 -530 60 -510
rect 100 -515 115 -495
rect 135 -515 160 -495
rect 100 -530 160 -515
rect 10 -555 60 -530
rect 110 -555 160 -530
rect 210 -555 260 -495
rect 390 -555 440 -495
rect 490 -555 540 -495
rect 590 -555 640 -495
rect 690 -555 740 -495
rect 870 -555 920 -495
rect 970 -555 1020 -495
rect 1070 -510 1120 -495
rect 1070 -530 1085 -510
rect 1105 -530 1120 -510
rect 1070 -555 1120 -530
rect 1560 -660 1605 -610
rect 2205 -660 2220 -610
rect 1560 -710 1580 -660
rect 1525 -725 1605 -710
rect 1525 -745 1540 -725
rect 1560 -745 1605 -725
rect 1525 -760 1605 -745
rect 2205 -760 2220 -710
rect 10 -880 60 -855
rect 110 -880 160 -855
rect 210 -880 260 -855
rect 390 -880 440 -855
rect 490 -880 540 -855
rect 590 -880 640 -855
rect 690 -880 740 -855
rect 870 -880 920 -855
rect 970 -880 1020 -855
rect 1070 -880 1120 -855
rect 865 -965 905 -955
rect 865 -985 875 -965
rect 895 -980 905 -965
rect 985 -965 1025 -955
rect 985 -980 995 -965
rect 895 -985 995 -980
rect 1015 -985 1025 -965
rect 865 -995 1025 -985
rect 485 -1025 525 -1015
rect 485 -1045 495 -1025
rect 515 -1040 525 -1025
rect 615 -1025 655 -1015
rect 1450 -1020 1500 -1010
rect 615 -1040 625 -1025
rect 515 -1045 625 -1040
rect 645 -1045 655 -1025
rect 485 -1055 655 -1045
rect 1340 -1030 1400 -1020
rect 1340 -1050 1350 -1030
rect 1370 -1050 1400 -1030
rect 1340 -1060 1400 -1050
rect 1350 -1075 1400 -1060
rect 1450 -1040 1460 -1020
rect 1480 -1040 1500 -1020
rect 1450 -1075 1500 -1040
rect 2260 -1020 2320 -1010
rect 2260 -1040 2290 -1020
rect 2310 -1040 2320 -1020
rect 2260 -1050 2320 -1040
rect 1550 -1075 1600 -1050
rect 1655 -1075 1705 -1050
rect 1755 -1075 1805 -1050
rect 1855 -1075 1905 -1050
rect 1955 -1075 2005 -1050
rect 2060 -1075 2110 -1050
rect 2160 -1075 2210 -1050
rect 2260 -1075 2310 -1050
rect 100 -1095 1020 -1080
rect 10 -1115 60 -1100
rect 10 -1135 25 -1115
rect 45 -1135 60 -1115
rect 100 -1115 115 -1095
rect 135 -1115 160 -1095
rect 100 -1130 160 -1115
rect 10 -1155 60 -1135
rect 110 -1155 160 -1130
rect 210 -1155 260 -1095
rect 390 -1155 440 -1095
rect 490 -1155 540 -1095
rect 590 -1155 640 -1095
rect 690 -1155 740 -1095
rect 870 -1155 920 -1095
rect 970 -1155 1020 -1095
rect 1070 -1115 1120 -1100
rect 1070 -1135 1085 -1115
rect 1105 -1135 1120 -1115
rect 1070 -1155 1120 -1135
rect 1350 -1390 1400 -1375
rect 1450 -1435 1500 -1375
rect 1550 -1435 1600 -1375
rect 1655 -1435 1705 -1375
rect 1755 -1435 1805 -1375
rect 1855 -1435 1905 -1375
rect 1955 -1435 2005 -1375
rect 2060 -1435 2110 -1375
rect 2160 -1435 2210 -1375
rect 2260 -1390 2310 -1375
rect 1450 -1450 2210 -1435
rect 10 -1480 60 -1455
rect 110 -1480 160 -1455
rect 210 -1480 260 -1455
rect 390 -1480 440 -1455
rect 490 -1480 540 -1455
rect 590 -1480 640 -1455
rect 690 -1480 740 -1455
rect 870 -1480 920 -1455
rect 970 -1480 1020 -1455
rect 1070 -1480 1120 -1455
rect 1740 -1490 1910 -1480
rect 1740 -1510 1750 -1490
rect 1770 -1495 1880 -1490
rect 1770 -1510 1780 -1495
rect 1740 -1520 1780 -1510
rect 1870 -1510 1880 -1495
rect 1900 -1510 1910 -1490
rect 1870 -1520 1910 -1510
<< polycont >>
rect 25 120 45 140
rect 125 135 145 155
rect 225 135 245 155
rect 325 135 345 155
rect 425 135 445 155
rect 525 135 545 155
rect 625 135 645 155
rect 725 135 745 155
rect 825 135 845 155
rect 925 120 945 140
rect 415 -285 435 -265
rect 675 -285 695 -265
rect 935 -285 955 -265
rect 1365 -345 1385 -325
rect 1455 -345 1475 -325
rect 2265 -345 2285 -325
rect 495 -425 515 -405
rect 615 -425 635 -405
rect 1455 -425 1475 -405
rect 1615 -425 1635 -405
rect 2015 -425 2035 -405
rect 2090 -415 2110 -395
rect 25 -530 45 -510
rect 115 -515 135 -495
rect 1085 -530 1105 -510
rect 1540 -745 1560 -725
rect 875 -985 895 -965
rect 995 -985 1015 -965
rect 495 -1045 515 -1025
rect 625 -1045 645 -1025
rect 1350 -1050 1370 -1030
rect 1460 -1040 1480 -1020
rect 2290 -1040 2310 -1020
rect 25 -1135 45 -1115
rect 115 -1115 135 -1095
rect 1085 -1135 1105 -1115
rect 1750 -1510 1770 -1490
rect 1880 -1510 1900 -1490
<< locali >>
rect 115 155 855 165
rect 15 140 55 150
rect 15 120 25 140
rect 45 120 55 140
rect 115 135 125 155
rect 145 135 225 155
rect 245 135 325 155
rect 345 135 425 155
rect 445 135 525 155
rect 545 135 625 155
rect 645 135 725 155
rect 745 135 825 155
rect 845 135 855 155
rect 115 125 855 135
rect 915 140 955 150
rect 15 110 55 120
rect 915 120 925 140
rect 945 120 955 140
rect 915 110 955 120
rect -85 80 5 90
rect -85 -190 -75 80
rect -55 -190 -25 80
rect -5 -190 5 80
rect -85 -200 5 -190
rect 65 80 105 90
rect 65 -190 75 80
rect 95 -190 105 80
rect 65 -395 105 -190
rect 165 80 205 90
rect 165 -190 175 80
rect 195 -190 205 80
rect 165 -200 205 -190
rect 265 80 305 90
rect 265 -190 275 80
rect 295 -190 305 80
rect 265 -255 305 -190
rect 365 80 405 90
rect 365 -190 375 80
rect 395 -190 405 80
rect 365 -200 405 -190
rect 465 80 505 90
rect 465 -190 475 80
rect 495 -190 505 80
rect 265 -265 445 -255
rect 265 -285 415 -265
rect 435 -285 445 -265
rect 265 -295 445 -285
rect 465 -395 505 -190
rect 565 80 605 90
rect 565 -190 575 80
rect 595 -190 605 80
rect 565 -200 605 -190
rect 665 80 705 90
rect 665 -190 675 80
rect 695 -190 705 80
rect 665 -255 705 -190
rect 765 80 805 90
rect 765 -190 775 80
rect 795 -190 805 80
rect 765 -200 805 -190
rect 865 80 905 90
rect 865 -190 875 80
rect 895 -190 905 80
rect 545 -265 705 -255
rect 545 -285 675 -265
rect 695 -285 705 -265
rect 545 -295 705 -285
rect 65 -405 525 -395
rect 65 -425 495 -405
rect 515 -425 525 -405
rect 65 -430 525 -425
rect 165 -435 525 -430
rect 105 -495 145 -485
rect 15 -510 55 -500
rect 15 -530 25 -510
rect 45 -530 55 -510
rect 105 -515 115 -495
rect 135 -515 145 -495
rect 105 -525 145 -515
rect 15 -540 55 -530
rect -85 -570 5 -560
rect -85 -840 -75 -570
rect -55 -840 -25 -570
rect -5 -840 5 -570
rect -85 -850 5 -840
rect 65 -570 105 -560
rect 65 -840 75 -570
rect 95 -840 105 -570
rect 65 -880 105 -840
rect 165 -570 205 -435
rect 545 -490 585 -295
rect 865 -395 905 -190
rect 965 80 1055 90
rect 965 -190 975 80
rect 995 -190 1025 80
rect 1045 -190 1055 80
rect 965 -200 1055 -190
rect 1195 20 2245 60
rect 1195 -255 1235 20
rect 925 -265 1235 -255
rect 925 -285 935 -265
rect 955 -285 1235 -265
rect 925 -295 1235 -285
rect 1255 -20 1345 -10
rect 1255 -290 1265 -20
rect 1285 -290 1315 -20
rect 1335 -290 1345 -20
rect 1255 -300 1345 -290
rect 1405 -20 1445 20
rect 1405 -290 1415 -20
rect 1435 -290 1445 -20
rect 1405 -295 1445 -290
rect 1505 -20 1545 -10
rect 1505 -290 1515 -20
rect 1535 -290 1545 -20
rect 1355 -325 1395 -315
rect 1355 -345 1365 -325
rect 1385 -345 1395 -325
rect 1355 -355 1395 -345
rect 1445 -325 1485 -315
rect 1445 -345 1455 -325
rect 1475 -345 1485 -325
rect 1445 -355 1485 -345
rect 605 -405 1485 -395
rect 605 -425 615 -405
rect 635 -425 1455 -405
rect 1475 -425 1485 -405
rect 605 -435 1485 -425
rect 445 -530 685 -490
rect 165 -840 175 -570
rect 195 -840 205 -570
rect 165 -850 205 -840
rect 265 -570 305 -560
rect 265 -840 275 -570
rect 295 -840 305 -570
rect 265 -880 305 -840
rect 65 -920 305 -880
rect 345 -570 385 -560
rect 345 -840 355 -570
rect 375 -840 385 -570
rect 345 -880 385 -840
rect 445 -570 485 -530
rect 445 -840 455 -570
rect 475 -840 485 -570
rect 445 -850 485 -840
rect 545 -570 585 -560
rect 545 -840 555 -570
rect 575 -840 585 -570
rect 545 -880 585 -840
rect 645 -570 685 -530
rect 645 -840 655 -570
rect 675 -840 685 -570
rect 645 -850 685 -840
rect 745 -570 785 -560
rect 745 -840 755 -570
rect 775 -840 785 -570
rect 745 -880 785 -840
rect 345 -920 785 -880
rect 825 -570 865 -560
rect 825 -840 835 -570
rect 855 -840 865 -570
rect 825 -880 865 -840
rect 925 -570 965 -435
rect 1505 -455 1545 -290
rect 1605 -20 1645 -10
rect 1605 -290 1615 -20
rect 1635 -290 1645 -20
rect 1605 -405 1645 -290
rect 1605 -425 1615 -405
rect 1635 -425 1645 -405
rect 1605 -435 1645 -425
rect 1705 -20 1745 -10
rect 1705 -290 1715 -20
rect 1735 -290 1745 -20
rect 1705 -455 1745 -290
rect 1805 -20 1845 20
rect 1805 -290 1815 -20
rect 1835 -290 1845 -20
rect 1805 -295 1845 -290
rect 1905 -20 1945 -10
rect 1905 -290 1915 -20
rect 1935 -290 1945 -20
rect 1905 -455 1945 -290
rect 2005 -20 2045 -10
rect 2005 -290 2015 -20
rect 2035 -290 2045 -20
rect 2005 -405 2045 -290
rect 2105 -20 2145 -10
rect 2105 -290 2115 -20
rect 2135 -290 2145 -20
rect 2105 -320 2145 -290
rect 2205 -20 2245 20
rect 2205 -290 2215 -20
rect 2235 -290 2245 -20
rect 2205 -295 2245 -290
rect 2305 -20 2395 -10
rect 2305 -290 2315 -20
rect 2335 -290 2365 -20
rect 2385 -290 2395 -20
rect 2305 -300 2395 -290
rect 2105 -360 2185 -320
rect 2255 -325 2295 -315
rect 2255 -345 2265 -325
rect 2285 -345 2295 -325
rect 2255 -355 2295 -345
rect 2005 -425 2015 -405
rect 2035 -425 2045 -405
rect 2080 -395 2120 -385
rect 2080 -415 2090 -395
rect 2110 -415 2120 -395
rect 2080 -425 2120 -415
rect 2005 -435 2045 -425
rect 2145 -455 2185 -360
rect 1505 -495 2260 -455
rect 1075 -510 1115 -500
rect 1075 -530 1085 -510
rect 1105 -530 1115 -510
rect 1075 -540 1115 -530
rect 925 -840 935 -570
rect 955 -840 965 -570
rect 925 -850 965 -840
rect 1025 -570 1065 -560
rect 1025 -840 1035 -570
rect 1055 -840 1065 -570
rect 1025 -880 1065 -840
rect 1125 -570 1215 -560
rect 2220 -565 2260 -495
rect 1125 -840 1135 -570
rect 1155 -840 1185 -570
rect 1205 -840 1215 -570
rect 1610 -575 2260 -565
rect 1610 -595 1620 -575
rect 2190 -595 2260 -575
rect 1610 -605 2260 -595
rect 1610 -675 2200 -665
rect 1610 -695 1620 -675
rect 2190 -695 2200 -675
rect 1610 -705 2200 -695
rect 1530 -725 1570 -715
rect 1530 -745 1540 -725
rect 1560 -745 1570 -725
rect 1530 -755 1570 -745
rect 2220 -765 2260 -605
rect 1610 -775 2260 -765
rect 1610 -795 1620 -775
rect 2190 -795 2260 -775
rect 1610 -805 2260 -795
rect 1125 -850 1215 -840
rect 825 -920 1065 -880
rect 165 -985 205 -920
rect 165 -1005 175 -985
rect 195 -1005 205 -985
rect 165 -1015 205 -1005
rect 545 -955 585 -920
rect 545 -965 905 -955
rect 545 -985 875 -965
rect 895 -985 905 -965
rect 545 -995 905 -985
rect 165 -1025 525 -1015
rect 165 -1045 495 -1025
rect 515 -1045 525 -1025
rect 165 -1055 525 -1045
rect 105 -1095 145 -1085
rect 15 -1115 55 -1105
rect 15 -1135 25 -1115
rect 45 -1135 55 -1115
rect 105 -1115 115 -1095
rect 135 -1115 145 -1095
rect 105 -1125 145 -1115
rect 15 -1145 55 -1135
rect -85 -1170 5 -1160
rect -85 -1440 -75 -1170
rect -55 -1440 -25 -1170
rect -5 -1440 5 -1170
rect -85 -1450 5 -1440
rect 65 -1170 105 -1160
rect 65 -1440 75 -1170
rect 95 -1440 105 -1170
rect 65 -1480 105 -1440
rect 165 -1170 205 -1055
rect 545 -1090 585 -995
rect 925 -1015 965 -920
rect 985 -965 1490 -955
rect 985 -985 995 -965
rect 1015 -985 1490 -965
rect 985 -995 1490 -985
rect 615 -1025 965 -1015
rect 1450 -1020 1490 -995
rect 615 -1045 625 -1025
rect 645 -1045 965 -1025
rect 615 -1055 965 -1045
rect 445 -1130 685 -1090
rect 165 -1440 175 -1170
rect 195 -1440 205 -1170
rect 165 -1450 205 -1440
rect 265 -1170 305 -1160
rect 265 -1440 275 -1170
rect 295 -1440 305 -1170
rect 265 -1480 305 -1440
rect 65 -1520 305 -1480
rect 345 -1170 385 -1160
rect 345 -1440 355 -1170
rect 375 -1440 385 -1170
rect 345 -1480 385 -1440
rect 445 -1170 485 -1130
rect 445 -1440 455 -1170
rect 475 -1440 485 -1170
rect 445 -1450 485 -1440
rect 545 -1170 585 -1160
rect 545 -1440 555 -1170
rect 575 -1440 585 -1170
rect 545 -1480 585 -1440
rect 645 -1170 685 -1130
rect 645 -1440 655 -1170
rect 675 -1440 685 -1170
rect 645 -1450 685 -1440
rect 745 -1170 785 -1160
rect 745 -1440 755 -1170
rect 775 -1440 785 -1170
rect 745 -1480 785 -1440
rect 345 -1520 785 -1480
rect 825 -1170 865 -1160
rect 825 -1440 835 -1170
rect 855 -1440 865 -1170
rect 825 -1480 865 -1440
rect 925 -1170 965 -1055
rect 1340 -1030 1380 -1020
rect 1340 -1050 1350 -1030
rect 1370 -1050 1380 -1030
rect 1450 -1040 1460 -1020
rect 1480 -1040 1490 -1020
rect 1450 -1050 1490 -1040
rect 2280 -1020 2320 -1010
rect 2280 -1040 2290 -1020
rect 2310 -1040 2320 -1020
rect 2280 -1050 2320 -1040
rect 1340 -1060 1380 -1050
rect 1255 -1090 1345 -1080
rect 1075 -1115 1115 -1105
rect 1075 -1135 1085 -1115
rect 1105 -1135 1115 -1115
rect 1075 -1145 1115 -1135
rect 925 -1440 935 -1170
rect 955 -1440 965 -1170
rect 925 -1450 965 -1440
rect 1025 -1170 1065 -1160
rect 1025 -1440 1035 -1170
rect 1055 -1440 1065 -1170
rect 1025 -1480 1065 -1440
rect 1125 -1170 1215 -1160
rect 1125 -1440 1135 -1170
rect 1155 -1440 1185 -1170
rect 1205 -1440 1215 -1170
rect 1255 -1360 1265 -1090
rect 1285 -1360 1315 -1090
rect 1335 -1360 1345 -1090
rect 1255 -1370 1345 -1360
rect 1405 -1090 1445 -1080
rect 1405 -1360 1415 -1090
rect 1435 -1360 1445 -1090
rect 1405 -1370 1445 -1360
rect 1505 -1090 1545 -1080
rect 1505 -1360 1515 -1090
rect 1535 -1360 1545 -1090
rect 1125 -1450 1215 -1440
rect 1505 -1480 1545 -1360
rect 1605 -1090 1650 -1080
rect 1605 -1360 1620 -1090
rect 1640 -1360 1650 -1090
rect 1605 -1370 1650 -1360
rect 1710 -1090 1750 -1080
rect 1710 -1360 1720 -1090
rect 1740 -1360 1750 -1090
rect 1710 -1400 1750 -1360
rect 1810 -1090 1850 -1080
rect 1810 -1360 1820 -1090
rect 1840 -1360 1850 -1090
rect 1810 -1370 1850 -1360
rect 1910 -1090 1950 -1080
rect 1910 -1360 1920 -1090
rect 1940 -1360 1950 -1090
rect 1910 -1400 1950 -1360
rect 2010 -1090 2055 -1080
rect 2010 -1360 2025 -1090
rect 2045 -1360 2055 -1090
rect 2010 -1370 2055 -1360
rect 2115 -1090 2155 -1080
rect 2115 -1360 2125 -1090
rect 2145 -1360 2155 -1090
rect 1710 -1440 1950 -1400
rect 825 -1490 1780 -1480
rect 825 -1510 1750 -1490
rect 1770 -1510 1780 -1490
rect 825 -1520 1780 -1510
rect 745 -1540 785 -1520
rect 1810 -1540 1850 -1440
rect 2115 -1480 2155 -1360
rect 2215 -1090 2255 -1080
rect 2215 -1360 2225 -1090
rect 2245 -1360 2255 -1090
rect 2215 -1370 2255 -1360
rect 2315 -1090 2405 -1080
rect 2315 -1360 2325 -1090
rect 2345 -1360 2375 -1090
rect 2395 -1360 2405 -1090
rect 2315 -1370 2405 -1360
rect 1870 -1490 2155 -1480
rect 1870 -1510 1880 -1490
rect 1900 -1510 2155 -1490
rect 1870 -1520 2155 -1510
rect 745 -1575 1850 -1540
<< viali >>
rect 25 120 45 140
rect 425 135 445 155
rect 925 120 945 140
rect -75 -190 -55 80
rect -25 -190 -5 80
rect 175 -190 195 80
rect 375 -190 395 80
rect 575 -190 595 80
rect 775 -190 795 80
rect 25 -530 45 -510
rect 115 -515 135 -495
rect -75 -840 -55 -570
rect -25 -840 -5 -570
rect 975 -190 995 80
rect 1025 -190 1045 80
rect 1265 -290 1285 -20
rect 1315 -290 1335 -20
rect 1455 -345 1475 -325
rect 2315 -290 2335 -20
rect 2365 -290 2385 -20
rect 2265 -345 2285 -325
rect 2090 -415 2110 -395
rect 1085 -530 1105 -510
rect 1135 -840 1155 -570
rect 1185 -840 1205 -570
rect 1620 -695 2190 -675
rect 175 -1005 195 -985
rect 25 -1135 45 -1115
rect 115 -1115 135 -1095
rect -75 -1365 -55 -1170
rect -75 -1440 -55 -1365
rect -25 -1440 -5 -1170
rect 1350 -1050 1370 -1030
rect 2290 -1040 2310 -1020
rect 1085 -1135 1105 -1115
rect 1135 -1440 1155 -1170
rect 1185 -1440 1205 -1170
rect 1265 -1360 1285 -1090
rect 1315 -1360 1335 -1090
rect 1415 -1360 1435 -1090
rect 1620 -1360 1640 -1090
rect 1820 -1360 1840 -1090
rect 2025 -1360 2045 -1090
rect 2225 -1360 2245 -1090
rect 2325 -1360 2345 -1090
rect 2375 -1360 2395 -1090
<< metal1 >>
rect 410 155 460 165
rect 15 140 55 150
rect 15 120 25 140
rect 45 120 55 140
rect 410 135 425 155
rect 445 135 460 155
rect 410 125 460 135
rect 915 140 955 150
rect 15 90 55 120
rect 915 120 925 140
rect 945 120 955 140
rect 915 90 955 120
rect -85 80 1055 90
rect -85 -190 -75 80
rect -55 -190 -25 80
rect -5 -190 175 80
rect 195 -190 375 80
rect 395 -190 575 80
rect 595 -190 775 80
rect 795 -190 975 80
rect 995 -190 1025 80
rect 1045 -190 1055 80
rect -85 -200 1055 -190
rect 1255 -20 2395 -10
rect 105 -495 145 -485
rect 10 -510 60 -495
rect 10 -530 25 -510
rect 45 -530 60 -510
rect 105 -515 115 -495
rect 135 -515 145 -495
rect 105 -525 145 -515
rect 10 -560 60 -530
rect 260 -560 870 -200
rect 1255 -290 1265 -20
rect 1285 -290 1315 -20
rect 1335 -290 2315 -20
rect 2335 -290 2365 -20
rect 2385 -290 2395 -20
rect 1255 -300 2395 -290
rect 1355 -355 1395 -300
rect 1445 -325 1485 -315
rect 1445 -345 1455 -325
rect 1475 -345 1485 -325
rect 1445 -355 1485 -345
rect 1075 -510 1115 -500
rect 1075 -530 1085 -510
rect 1105 -530 1115 -510
rect 1075 -560 1115 -530
rect -85 -570 1215 -560
rect -85 -840 -75 -570
rect -55 -840 -25 -570
rect -5 -840 1135 -570
rect 1155 -840 1185 -570
rect 1205 -840 1215 -570
rect 1600 -665 2050 -300
rect 2255 -325 2295 -300
rect 2255 -345 2265 -325
rect 2285 -345 2295 -325
rect 2255 -355 2295 -345
rect 2080 -395 2120 -385
rect 2080 -415 2090 -395
rect 2110 -415 2120 -395
rect 2080 -425 2120 -415
rect 1600 -675 2200 -665
rect 1600 -695 1620 -675
rect 2190 -695 2200 -675
rect 1600 -705 2200 -695
rect 1530 -755 1570 -715
rect -85 -850 1215 -840
rect -85 -855 1050 -850
rect 165 -985 205 -975
rect 165 -1005 175 -985
rect 195 -1005 205 -985
rect 165 -1015 205 -1005
rect 1075 -1030 1395 -1020
rect 1075 -1050 1350 -1030
rect 1370 -1050 1395 -1030
rect 1075 -1075 1395 -1050
rect 1600 -1075 2050 -705
rect 2265 -1020 2320 -1010
rect 2265 -1040 2290 -1020
rect 2310 -1040 2320 -1020
rect 2265 -1050 2320 -1040
rect 2265 -1075 2310 -1050
rect 1075 -1080 2310 -1075
rect 105 -1095 145 -1085
rect 15 -1115 55 -1105
rect 15 -1135 25 -1115
rect 45 -1135 55 -1115
rect 105 -1115 115 -1095
rect 135 -1115 145 -1095
rect 105 -1125 145 -1115
rect 1075 -1090 2405 -1080
rect 1075 -1115 1265 -1090
rect 15 -1160 55 -1135
rect 1075 -1135 1085 -1115
rect 1105 -1135 1265 -1115
rect 1075 -1160 1265 -1135
rect -85 -1170 1265 -1160
rect -85 -1440 -75 -1170
rect -55 -1440 -25 -1170
rect -5 -1440 1135 -1170
rect 1155 -1440 1185 -1170
rect 1205 -1360 1265 -1170
rect 1285 -1360 1315 -1090
rect 1335 -1360 1415 -1090
rect 1435 -1360 1620 -1090
rect 1640 -1360 1820 -1090
rect 1840 -1360 2025 -1090
rect 2045 -1360 2225 -1090
rect 2245 -1360 2325 -1090
rect 2345 -1360 2375 -1090
rect 2395 -1360 2405 -1090
rect 1205 -1370 2405 -1360
rect 1205 -1440 1395 -1370
rect -85 -1450 1395 -1440
<< labels >>
rlabel metal1 -85 -1305 -85 -1305 7 VN
port 2 w
rlabel metal1 410 145 410 145 7 VBP
port 3 w
rlabel metal1 105 -505 105 -505 3 VCP
port 4 e
rlabel metal1 105 -1105 105 -1105 3 VCN
port 5 e
rlabel metal1 1530 -735 1530 -735 7 VBN
port 8 w
rlabel metal1 165 -995 165 -995 7 VOUT
port 9 w
rlabel metal1 -85 -55 -85 -55 7 VP
port 1 w
rlabel metal1 1445 -335 1445 -335 3 V1
port 6 e
rlabel metal1 2080 -405 2080 -405 7 V2
port 7 w
<< end >>
