* NGSPICE file created from top_differential_amplifier.ext - technology: sky130A

.subckt bias_generator VP VN VBP VBN VCN VCP
X0 a_2450_n4910# VCN VCN VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X1 VN VBN VCP VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X2 VBP VBP VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X3 a_5640_n2240# a_5740_n2350# a_5740_n2350# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X4 VBP VBP VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X5 a_5640_n2240# VCP VCP VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X6 VP a_5740_n2350# a_5640_n2240# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X7 a_3650_n2110# VBP a_2550_n4950# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X8 VCN VBP VP VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X9 a_2550_n4950# a_2550_n4950# a_2450_n4910# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X10 a_7440_n4910# VBN a_7240_n4910# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X11 a_2650_n2110# VBP VP VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X12 a_2450_n4910# a_2550_n4950# a_2550_n4950# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X13 VCP VN VN VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.4 ps=24.9 w=12 l=0.5
X14 a_6440_n4910# VBN a_6240_n4910# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X15 VCN VN VN VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=0.5
X16 a_5640_n2240# a_5740_n2350# a_5740_n2350# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X17 a_5740_n2350# a_5740_n2350# a_5640_n2240# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X18 VBN VBP VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X19 VP VBP a_4250_n2110# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X20 VCP VP VP VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=5.4 ps=24.9 w=12 l=0.5
X21 a_2550_n4950# VBP a_3250_n2110# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X22 a_7240_n4910# VBN a_7040_n4910# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X23 VP VBP VCN VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X24 a_6240_n4910# VBN a_6040_n4910# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X25 VP VBP VBN VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X26 a_5740_n2350# a_5740_n2350# a_5640_n2240# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X27 a_5640_n2240# a_5740_n2350# a_5740_n2350# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X28 a_2550_n4950# a_2550_n4950# a_2450_n4910# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X29 a_2450_n4910# a_2550_n4950# a_2550_n4950# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X30 VP VBP VBN VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X31 a_4250_n2110# VBP a_4050_n2110# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X32 a_3250_n2110# VBP a_3050_n2110# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X33 VCN VP VP VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=0.5
X34 VP VP VBN VP sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=0.75 ps=3.5 w=3 l=0.5
X35 a_2550_n4950# a_2550_n4950# a_2450_n4910# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X36 VN VN VCN VN sky130_fd_pr__nfet_01v8 ad=5.4 pd=24.9 as=3 ps=12.5 w=12 l=0.5
X37 a_7040_n4910# VBN a_6840_n4910# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X38 VN VN VCP VN sky130_fd_pr__nfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=0.5
X39 a_2450_n4910# a_2550_n4950# a_2550_n4950# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X40 a_6040_n4910# VBN a_5840_n4910# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X41 VP VBP VBP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X42 VP VBP VBP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X43 VP VP VCP VP sky130_fd_pr__pfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=0.5
X44 a_5740_n2350# a_5740_n2350# a_5640_n2240# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X45 a_5640_n2240# a_5740_n2350# a_5740_n2350# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X46 VCP VBN VN VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X47 a_3050_n2110# VBP a_2850_n2110# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X48 a_4050_n2110# VBP a_3850_n2110# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X49 VN VBN VBN VN sky130_fd_pr__nfet_01v8 ad=6 pd=25 as=6 ps=25 w=12 l=0.5
X50 a_2450_n4910# a_2550_n4950# VN VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X51 VCN VCN a_2450_n4910# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X52 a_6840_n4910# VBN a_5740_n2350# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X53 VBN VBP VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X54 a_2550_n4950# a_2550_n4950# a_2450_n4910# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X55 a_5840_n4910# VBN VN VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X56 VBN VP VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.5 ps=7 w=3 l=0.5
X57 VCP VCP a_5640_n2240# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X58 a_5640_n2240# a_5740_n2350# VP VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X59 VP VP VCN VP sky130_fd_pr__pfet_01v8 ad=5.4 pd=24.9 as=3 ps=12.5 w=12 l=0.5
X60 a_5740_n2350# a_5740_n2350# a_5640_n2240# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X61 a_2450_n4910# a_2550_n4950# a_2550_n4950# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X62 VN VBN a_7440_n4910# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X63 a_2850_n2110# VBP a_2650_n2110# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X64 a_3850_n2110# VBP a_3650_n2110# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X65 VN a_2550_n4950# a_2450_n4910# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X66 a_5740_n2350# VBN a_6440_n4910# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
.ends

.subckt folded_cascode_differential_amplifier VP VN VBP VCP VCN V1 V2 VBN VOUT
X0 VN VN a_520_n410# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=0.5
X1 VOUT VP VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.5 ps=7 w=3 l=0.5
X2 a_520_n410# VCP a_680_n1710# VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X3 VOUT VCN a_120_n2910# VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X4 a_680_n2910# a_680_n1710# VN VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X5 a_120_n410# V2 a_3000_n610# VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X6 VN VBN a_3000_n610# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X7 a_520_n410# V1 a_3000_n610# VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X8 a_680_n1710# VCN a_680_n2910# VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.5 ps=7 w=3 l=0.5
X9 a_120_n410# V2 a_3000_n610# VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X10 a_120_n2910# a_680_n1710# VN VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X11 VN a_680_n1710# a_120_n2910# VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X12 a_3000_n610# V1 a_520_n410# VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X13 VN a_680_n1710# a_680_n2910# VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X14 VOUT VCP a_120_n410# VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X15 VP VBP a_120_n410# VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X16 VOUT VCP a_120_n410# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=0.5
X17 VP VBP a_520_n410# VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X18 VP VBP a_120_n410# VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X19 VN VN VN VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=19.8 ps=90.2 w=3 l=0.5
X20 a_120_n2910# a_680_n1710# VN VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.825 ps=3.55 w=3 l=0.5
X21 VP VBP a_520_n410# VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X22 VP VP a_120_n410# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=0.5
X23 a_680_n1710# VCP a_520_n410# VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X24 a_680_n2910# VCN a_680_n1710# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=0.5
X25 a_680_n2910# a_680_n1710# VN VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.825 ps=3.55 w=3 l=0.5
X26 a_120_n410# VP VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.5 ps=7 w=3 l=0.5
X27 a_120_n410# VCP VOUT VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.5 ps=7 w=3 l=0.5
X28 a_120_n410# VCP VOUT VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X29 a_520_n410# V1 a_3000_n610# VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X30 VN VN a_120_n2910# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=0.5
X31 a_680_n1710# VCN a_680_n2910# VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X32 a_3000_n610# V2 a_120_n410# VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X33 a_520_n410# VCP a_680_n1710# VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.5 ps=7 w=3 l=0.5
X34 a_120_n2910# VN VN VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.5 ps=7 w=3 l=0.5
X35 a_3000_n610# V1 a_520_n410# VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X36 a_520_n410# VN VN VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.5 ps=7 w=3 l=0.5
X37 a_3000_n610# VBN VN VN sky130_fd_pr__nfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X38 a_120_n2910# VCN VOUT VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X39 a_520_n410# VBP VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X40 a_120_n410# VBP VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X41 a_520_n410# VBP VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X42 a_680_n1710# VCP a_520_n410# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=0.5
X43 a_120_n2910# VCN VOUT VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=0.5
X44 a_120_n410# VBP VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X45 VN a_680_n1710# a_120_n2910# VN sky130_fd_pr__nfet_01v8 ad=0.825 pd=3.55 as=0.75 ps=3.5 w=3 l=0.5
X46 VN a_680_n1710# a_680_n2910# VN sky130_fd_pr__nfet_01v8 ad=0.825 pd=3.55 as=0.75 ps=3.5 w=3 l=0.5
X47 a_680_n2910# VCN a_680_n1710# VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X48 VP VP VOUT VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=0.5
X49 a_3000_n610# V2 a_120_n410# VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X50 VOUT VCN a_120_n2910# VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.5 ps=7 w=3 l=0.5
X51 VN VN VN VN sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0 ps=0 w=3 l=0.5
.ends


* Top level circuit top_differential_amplifier

Xbias_generator_0 VP VN IB bias_generator_0/VBN bias_generator_0/VCN bias_generator_0/VCP
+ bias_generator
Xfolded_cascode_differential_amplifier_0 VP VN IB bias_generator_0/VCP bias_generator_0/VCN
+ V1 V2 bias_generator_0/VBN VOUT folded_cascode_differential_amplifier
X0 VP IB IB VP sky130_fd_pr__pfet_01v8 ad=6 pd=25 as=6 ps=25 w=12 l=0.5
.end

