magic
tech sky130A
timestamp 1697385496
<< locali >>
rect -5 1870 35 1910
rect 3370 1425 3410 1465
rect 245 70 285 110
rect 575 0 615 40
<< metal1 >>
rect 55 2775 95 2815
rect 345 1275 385 1315
use bias_generator  bias_generator_0
timestamp 1697384475
transform 1 0 -555 0 1 2675
box 550 -2735 4140 205
<< labels >>
rlabel locali 245 90 245 90 7 VBN
rlabel locali 575 20 575 20 7 VCN
rlabel metal1 365 1315 365 1315 1 VN
rlabel locali -5 1890 -5 1890 7 VBP
rlabel metal1 55 2795 55 2795 7 VP
rlabel locali 3410 1445 3410 1445 3 VCP
<< end >>
