magic
tech sky130A
timestamp 1697311719
<< nmos >>
rect 10 -205 60 95
rect 110 -205 160 95
rect 210 -205 260 95
rect 310 -205 360 95
rect 410 -205 460 95
rect 510 -205 560 95
rect 610 -205 660 95
rect 710 -205 760 95
rect 810 -205 860 95
rect 910 -205 960 95
<< ndiff >>
rect -40 80 10 95
rect -40 -190 -25 80
rect -5 -190 10 80
rect -40 -205 10 -190
rect 60 80 110 95
rect 60 -190 75 80
rect 95 -190 110 80
rect 60 -205 110 -190
rect 160 80 210 95
rect 160 -190 175 80
rect 195 -190 210 80
rect 160 -205 210 -190
rect 260 80 310 95
rect 260 -190 275 80
rect 295 -190 310 80
rect 260 -205 310 -190
rect 360 80 410 95
rect 360 -190 375 80
rect 395 -190 410 80
rect 360 -205 410 -190
rect 460 80 510 95
rect 460 -190 475 80
rect 495 -190 510 80
rect 460 -205 510 -190
rect 560 80 610 95
rect 560 -190 575 80
rect 595 -190 610 80
rect 560 -205 610 -190
rect 660 80 710 95
rect 660 -190 675 80
rect 695 -190 710 80
rect 660 -205 710 -190
rect 760 80 810 95
rect 760 -190 775 80
rect 795 -190 810 80
rect 760 -205 810 -190
rect 860 80 910 95
rect 860 -190 875 80
rect 895 -190 910 80
rect 860 -205 910 -190
rect 960 80 1010 95
rect 960 -190 975 80
rect 995 -190 1010 80
rect 960 -205 1010 -190
<< ndiffc >>
rect -25 -190 -5 80
rect 75 -190 95 80
rect 175 -190 195 80
rect 275 -190 295 80
rect 375 -190 395 80
rect 475 -190 495 80
rect 575 -190 595 80
rect 675 -190 695 80
rect 775 -190 795 80
rect 875 -190 895 80
rect 975 -190 995 80
<< psubdiff >>
rect -90 80 -40 95
rect -90 -190 -75 80
rect -55 -190 -40 80
rect -90 -205 -40 -190
rect 1010 80 1060 95
rect 1010 -190 1025 80
rect 1045 -190 1060 80
rect 1010 -205 1060 -190
<< psubdiffcont >>
rect -75 -190 -55 80
rect 1025 -190 1045 80
<< poly >>
rect 10 155 60 170
rect 10 135 25 155
rect 45 135 60 155
rect 10 95 60 135
rect 110 155 160 170
rect 110 135 125 155
rect 145 135 160 155
rect 110 95 160 135
rect 210 155 260 170
rect 210 135 225 155
rect 245 135 260 155
rect 210 95 260 135
rect 310 155 360 170
rect 310 135 325 155
rect 345 135 360 155
rect 310 95 360 135
rect 410 155 460 170
rect 410 135 425 155
rect 445 135 460 155
rect 410 95 460 135
rect 510 155 560 170
rect 510 135 525 155
rect 545 135 560 155
rect 510 95 560 135
rect 610 155 660 170
rect 610 135 625 155
rect 645 135 660 155
rect 610 95 660 135
rect 710 155 760 170
rect 710 135 725 155
rect 745 135 760 155
rect 710 95 760 135
rect 810 155 860 170
rect 810 135 825 155
rect 845 135 860 155
rect 810 95 860 135
rect 910 155 960 170
rect 910 135 925 155
rect 945 135 960 155
rect 910 95 960 135
rect 10 -230 60 -205
rect 110 -230 160 -205
rect 210 -230 260 -205
rect 310 -230 360 -205
rect 410 -230 460 -205
rect 510 -230 560 -205
rect 610 -230 660 -205
rect 710 -230 760 -205
rect 810 -230 860 -205
rect 910 -230 960 -205
<< polycont >>
rect 25 135 45 155
rect 125 135 145 155
rect 225 135 245 155
rect 325 135 345 155
rect 425 135 445 155
rect 525 135 545 155
rect 625 135 645 155
rect 725 135 745 155
rect 825 135 845 155
rect 925 135 945 155
<< locali >>
rect 15 155 55 165
rect 15 135 25 155
rect 45 135 55 155
rect 15 125 55 135
rect 115 155 855 165
rect 115 135 125 155
rect 145 135 225 155
rect 245 135 325 155
rect 345 135 425 155
rect 445 135 525 155
rect 545 135 625 155
rect 645 135 725 155
rect 745 135 825 155
rect 845 135 855 155
rect 115 125 855 135
rect 915 155 955 165
rect 915 135 925 155
rect 945 135 955 155
rect 915 125 955 135
rect -85 80 5 90
rect -85 -190 -75 80
rect -55 -190 -25 80
rect -5 -190 5 80
rect -85 -200 5 -190
rect 65 80 105 90
rect 65 -190 75 80
rect 95 -190 105 80
rect 65 -200 105 -190
rect 165 80 205 90
rect 165 -190 175 80
rect 195 -190 205 80
rect 165 -200 205 -190
rect 265 80 305 90
rect 265 -190 275 80
rect 295 -190 305 80
rect 265 -200 305 -190
rect 365 80 405 90
rect 365 -190 375 80
rect 395 -190 405 80
rect 365 -200 405 -190
rect 465 80 505 90
rect 465 -190 475 80
rect 495 -190 505 80
rect 465 -200 505 -190
rect 565 80 605 90
rect 565 -190 575 80
rect 595 -190 605 80
rect 565 -200 605 -190
rect 665 80 705 90
rect 665 -190 675 80
rect 695 -190 705 80
rect 665 -200 705 -190
rect 765 80 805 90
rect 765 -190 775 80
rect 795 -190 805 80
rect 765 -200 805 -190
rect 865 80 905 90
rect 865 -190 875 80
rect 895 -190 905 80
rect 865 -200 905 -190
rect 965 80 1055 90
rect 965 -190 975 80
rect 995 -190 1025 80
rect 1045 -190 1055 80
rect 965 -200 1055 -190
<< viali >>
rect -75 -190 -55 80
rect -25 -190 -5 80
rect 175 -190 195 80
rect 375 -190 395 80
rect 575 -190 595 80
rect 775 -190 795 80
rect 975 -190 995 80
rect 1025 -190 1045 80
<< metal1 >>
rect -85 80 1055 90
rect -85 -190 -75 80
rect -55 -190 -25 80
rect -5 -190 175 80
rect 195 -190 375 80
rect 395 -190 575 80
rect 595 -190 775 80
rect 795 -190 975 80
rect 995 -190 1025 80
rect 1045 -190 1055 80
rect -85 -200 1055 -190
<< end >>
