magic
tech sky130A
timestamp 1695762812
use crsl_d_flip_flop  crsl_d_flip_flop_0
timestamp 1695762812
transform 1 0 80 0 1 1510
box -85 -1545 230 545
<< end >>
