magic
tech sky130A
timestamp 1695699366
<< error_p >>
rect 800 -525 836 -524
<< nwell >>
rect 85 -405 470 445
<< nmos >>
rect 645 495 745 510
rect 645 430 745 445
rect 645 285 745 300
rect 645 220 745 235
rect 645 15 745 30
rect 250 -540 265 -440
rect 250 -690 265 -590
rect 645 -130 745 -115
rect 645 -275 745 -260
rect 645 -680 745 -665
rect 185 -795 315 -780
rect 210 -1070 310 -1055
rect 210 -1135 310 -1120
rect 210 -1280 310 -1265
rect 210 -1345 310 -1330
rect 645 -825 745 -810
rect 645 -970 745 -955
rect 645 -1115 745 -1100
rect 645 -1180 745 -1165
rect 645 -1365 745 -1350
rect 645 -1430 745 -1415
<< pmos >>
rect 210 355 310 370
rect 210 290 310 305
rect 210 140 310 155
rect 210 75 310 90
rect 250 -105 265 -5
rect 250 -235 265 -135
rect 250 -385 265 -285
<< ndiff >>
rect 645 545 745 560
rect 645 525 660 545
rect 730 525 745 545
rect 645 510 745 525
rect 645 480 745 495
rect 645 460 660 480
rect 730 460 745 480
rect 645 445 745 460
rect 645 415 745 430
rect 645 395 660 415
rect 730 395 745 415
rect 645 380 745 395
rect 645 335 745 350
rect 645 315 660 335
rect 730 315 745 335
rect 645 300 745 315
rect 645 270 745 285
rect 645 250 660 270
rect 730 250 745 270
rect 645 235 745 250
rect 645 205 745 220
rect 645 185 660 205
rect 730 185 745 205
rect 645 170 745 185
rect 645 65 745 80
rect 645 45 660 65
rect 730 45 745 65
rect 645 30 745 45
rect 645 0 745 15
rect 645 -20 660 0
rect 730 -20 745 0
rect 200 -455 250 -440
rect 200 -525 215 -455
rect 235 -525 250 -455
rect 200 -540 250 -525
rect 265 -455 315 -440
rect 265 -525 280 -455
rect 300 -525 315 -455
rect 265 -540 315 -525
rect 200 -605 250 -590
rect 200 -675 215 -605
rect 235 -675 250 -605
rect 200 -690 250 -675
rect 265 -605 315 -590
rect 265 -675 280 -605
rect 300 -675 315 -605
rect 265 -690 315 -675
rect 645 -35 745 -20
rect 645 -80 745 -65
rect 645 -100 660 -80
rect 730 -100 745 -80
rect 645 -115 745 -100
rect 645 -145 745 -130
rect 645 -165 660 -145
rect 730 -165 745 -145
rect 645 -180 745 -165
rect 645 -225 745 -210
rect 645 -245 660 -225
rect 730 -245 745 -225
rect 645 -260 745 -245
rect 645 -290 745 -275
rect 645 -310 660 -290
rect 730 -310 745 -290
rect 645 -325 745 -310
rect 645 -630 745 -615
rect 645 -650 660 -630
rect 730 -650 745 -630
rect 645 -665 745 -650
rect 645 -695 745 -680
rect 185 -745 315 -730
rect 185 -765 200 -745
rect 300 -765 315 -745
rect 185 -780 315 -765
rect 185 -810 315 -795
rect 185 -830 200 -810
rect 300 -830 315 -810
rect 185 -845 315 -830
rect 210 -1020 310 -1005
rect 210 -1040 225 -1020
rect 295 -1040 310 -1020
rect 210 -1055 310 -1040
rect 210 -1085 310 -1070
rect 210 -1105 225 -1085
rect 295 -1105 310 -1085
rect 210 -1120 310 -1105
rect 210 -1150 310 -1135
rect 210 -1170 225 -1150
rect 295 -1170 310 -1150
rect 210 -1185 310 -1170
rect 210 -1230 310 -1215
rect 210 -1250 225 -1230
rect 295 -1250 310 -1230
rect 210 -1265 310 -1250
rect 210 -1295 310 -1280
rect 210 -1315 225 -1295
rect 295 -1315 310 -1295
rect 210 -1330 310 -1315
rect 210 -1360 310 -1345
rect 210 -1380 225 -1360
rect 295 -1380 310 -1360
rect 210 -1395 310 -1380
rect 645 -715 660 -695
rect 730 -715 745 -695
rect 645 -730 745 -715
rect 645 -775 745 -760
rect 645 -795 660 -775
rect 730 -795 745 -775
rect 645 -810 745 -795
rect 645 -840 745 -825
rect 645 -860 660 -840
rect 730 -860 745 -840
rect 645 -875 745 -860
rect 645 -920 745 -905
rect 645 -940 660 -920
rect 730 -940 745 -920
rect 645 -955 745 -940
rect 645 -985 745 -970
rect 645 -1005 660 -985
rect 730 -1005 745 -985
rect 645 -1020 745 -1005
rect 645 -1065 745 -1050
rect 645 -1085 660 -1065
rect 730 -1085 745 -1065
rect 645 -1100 745 -1085
rect 645 -1130 745 -1115
rect 645 -1150 660 -1130
rect 730 -1150 745 -1130
rect 645 -1165 745 -1150
rect 645 -1195 745 -1180
rect 645 -1215 660 -1195
rect 730 -1215 745 -1195
rect 645 -1230 745 -1215
rect 645 -1315 745 -1300
rect 645 -1335 660 -1315
rect 730 -1335 745 -1315
rect 645 -1350 745 -1335
rect 645 -1380 745 -1365
rect 645 -1400 660 -1380
rect 730 -1400 745 -1380
rect 645 -1415 745 -1400
rect 645 -1445 745 -1430
rect 645 -1465 660 -1445
rect 730 -1465 745 -1445
rect 645 -1480 745 -1465
<< pdiff >>
rect 210 405 310 420
rect 210 385 225 405
rect 295 385 310 405
rect 210 370 310 385
rect 210 340 310 355
rect 210 320 225 340
rect 295 320 310 340
rect 210 305 310 320
rect 210 275 310 290
rect 210 255 225 275
rect 295 255 310 275
rect 210 240 310 255
rect 210 190 310 205
rect 210 170 225 190
rect 295 170 310 190
rect 210 155 310 170
rect 210 125 310 140
rect 210 105 225 125
rect 295 105 310 125
rect 210 90 310 105
rect 210 60 310 75
rect 210 40 225 60
rect 295 40 310 60
rect 210 25 310 40
rect 200 -20 250 -5
rect 200 -90 215 -20
rect 235 -90 250 -20
rect 200 -105 250 -90
rect 265 -20 315 -5
rect 265 -90 280 -20
rect 300 -90 315 -20
rect 265 -105 315 -90
rect 200 -150 250 -135
rect 200 -220 215 -150
rect 235 -220 250 -150
rect 200 -235 250 -220
rect 265 -150 315 -135
rect 265 -220 280 -150
rect 300 -220 315 -150
rect 265 -235 315 -220
rect 200 -300 250 -285
rect 200 -370 215 -300
rect 235 -370 250 -300
rect 200 -385 250 -370
rect 265 -300 315 -285
rect 265 -370 280 -300
rect 300 -370 315 -300
rect 265 -385 315 -370
<< ndiffc >>
rect 660 525 730 545
rect 660 460 730 480
rect 660 395 730 415
rect 660 315 730 335
rect 660 250 730 270
rect 660 185 730 205
rect 660 45 730 65
rect 660 -20 730 0
rect 215 -525 235 -455
rect 280 -525 300 -455
rect 215 -675 235 -605
rect 280 -675 300 -605
rect 660 -100 730 -80
rect 660 -165 730 -145
rect 660 -245 730 -225
rect 660 -310 730 -290
rect 660 -650 730 -630
rect 200 -765 300 -745
rect 200 -830 300 -810
rect 225 -1040 295 -1020
rect 225 -1105 295 -1085
rect 225 -1170 295 -1150
rect 225 -1250 295 -1230
rect 225 -1315 295 -1295
rect 225 -1380 295 -1360
rect 660 -715 730 -695
rect 660 -795 730 -775
rect 660 -860 730 -840
rect 660 -940 730 -920
rect 660 -1005 730 -985
rect 660 -1085 730 -1065
rect 660 -1150 730 -1130
rect 660 -1215 730 -1195
rect 660 -1335 730 -1315
rect 660 -1400 730 -1380
rect 660 -1465 730 -1445
<< pdiffc >>
rect 225 385 295 405
rect 225 320 295 340
rect 225 255 295 275
rect 225 170 295 190
rect 225 105 295 125
rect 225 40 295 60
rect 215 -90 235 -20
rect 280 -90 300 -20
rect 215 -220 235 -150
rect 280 -220 300 -150
rect 215 -370 235 -300
rect 280 -370 300 -300
<< psubdiff >>
rect 545 315 595 415
rect 625 -545 675 -445
rect 240 -890 290 -875
rect 240 -960 255 -890
rect 275 -960 290 -890
rect 240 -975 290 -960
<< nsubdiff >>
rect 380 410 430 425
rect 380 340 395 410
rect 415 340 430 410
rect 380 325 430 340
<< psubdiffcont >>
rect 255 -960 275 -890
<< nsubdiffcont >>
rect 395 340 415 410
<< poly >>
rect 590 500 645 510
rect 590 480 600 500
rect 620 495 645 500
rect 745 495 760 510
rect 620 480 630 495
rect 590 470 630 480
rect 630 430 645 445
rect 745 435 800 445
rect 745 430 770 435
rect 195 355 210 370
rect 310 360 365 370
rect 310 355 335 360
rect 115 320 155 330
rect 115 300 125 320
rect 145 305 155 320
rect 325 340 335 355
rect 355 340 365 360
rect 325 330 365 340
rect 760 415 770 430
rect 790 415 800 435
rect 760 405 800 415
rect 760 355 800 365
rect 760 335 770 355
rect 790 335 800 355
rect 760 325 800 335
rect 145 300 210 305
rect 115 290 210 300
rect 310 290 405 305
rect 155 220 340 230
rect 155 215 365 220
rect 155 90 170 215
rect 325 210 365 215
rect 325 190 335 210
rect 355 190 365 210
rect 325 180 365 190
rect 195 140 210 155
rect 310 145 365 155
rect 310 140 335 145
rect 325 125 335 140
rect 355 125 365 145
rect 325 115 365 125
rect 155 75 210 90
rect 310 75 325 90
rect 105 -105 145 -95
rect 105 -125 115 -105
rect 135 -125 145 -105
rect 105 -135 145 -125
rect 105 -355 120 -135
rect 170 -230 185 75
rect 250 -5 265 10
rect 250 -135 265 -105
rect 145 -240 185 -230
rect 390 -180 405 290
rect 550 290 645 300
rect 550 270 560 290
rect 580 285 645 290
rect 745 285 760 300
rect 580 270 590 285
rect 550 260 590 270
rect 785 235 800 325
rect 630 220 645 235
rect 745 220 800 235
rect 590 185 630 195
rect 590 165 600 185
rect 620 165 630 185
rect 590 155 630 165
rect 615 95 630 155
rect 590 85 630 95
rect 590 65 600 85
rect 620 65 630 85
rect 590 55 630 65
rect 785 70 800 220
rect 785 55 815 70
rect 630 15 645 30
rect 745 15 775 30
rect 550 5 590 15
rect 550 -15 560 5
rect 580 -15 590 5
rect 550 -25 590 -15
rect 390 -195 410 -180
rect 145 -260 155 -240
rect 175 -260 185 -240
rect 145 -270 185 -260
rect 105 -365 145 -355
rect 105 -385 115 -365
rect 135 -385 145 -365
rect 105 -395 145 -385
rect 170 -445 185 -270
rect 250 -285 265 -235
rect 330 -240 370 -230
rect 330 -260 340 -240
rect 360 -260 370 -240
rect 330 -270 370 -260
rect 250 -440 265 -385
rect 145 -455 185 -445
rect 145 -475 155 -455
rect 175 -475 185 -455
rect 145 -485 185 -475
rect 170 -700 185 -485
rect 250 -590 265 -540
rect 335 -545 350 -270
rect 395 -280 410 -195
rect 390 -295 410 -280
rect 390 -330 405 -295
rect 390 -340 430 -330
rect 390 -360 400 -340
rect 420 -360 430 -340
rect 390 -370 430 -360
rect 325 -555 365 -545
rect 325 -575 335 -555
rect 355 -575 365 -555
rect 325 -585 365 -575
rect 550 -665 565 -25
rect 590 -60 630 -50
rect 590 -80 600 -60
rect 620 -80 630 -60
rect 590 -90 630 -80
rect 590 -600 605 -90
rect 760 -115 775 15
rect 800 -5 815 55
rect 800 -15 840 -5
rect 800 -35 810 -15
rect 830 -35 840 -15
rect 800 -45 840 -35
rect 630 -130 645 -115
rect 745 -130 775 -115
rect 760 -260 775 -130
rect 800 -185 840 -175
rect 800 -205 810 -185
rect 830 -205 840 -185
rect 800 -215 840 -205
rect 630 -275 645 -260
rect 745 -275 775 -260
rect 760 -340 775 -275
rect 675 -350 775 -340
rect 675 -370 685 -350
rect 705 -355 775 -350
rect 705 -370 715 -355
rect 675 -380 715 -370
rect 700 -585 715 -380
rect 740 -390 780 -380
rect 740 -410 750 -390
rect 770 -410 780 -390
rect 740 -420 780 -410
rect 760 -545 775 -420
rect 825 -485 840 -215
rect 800 -495 840 -485
rect 800 -515 810 -495
rect 830 -515 840 -495
rect 800 -525 840 -515
rect 760 -560 815 -545
rect 700 -600 775 -585
rect 590 -610 630 -600
rect 590 -630 600 -610
rect 620 -630 630 -610
rect 590 -640 630 -630
rect 760 -665 775 -600
rect 550 -675 590 -665
rect 130 -715 185 -700
rect 250 -705 265 -690
rect 550 -695 560 -675
rect 580 -695 590 -675
rect 630 -680 645 -665
rect 745 -680 775 -665
rect 550 -705 590 -695
rect 130 -1095 145 -715
rect 250 -720 345 -705
rect 330 -780 345 -720
rect 170 -795 185 -780
rect 315 -795 345 -780
rect 330 -910 345 -795
rect 330 -925 450 -910
rect 195 -1070 210 -1055
rect 310 -1070 365 -1055
rect 130 -1105 195 -1095
rect 130 -1110 165 -1105
rect 155 -1125 165 -1110
rect 185 -1120 195 -1105
rect 185 -1125 210 -1120
rect 155 -1135 210 -1125
rect 310 -1135 325 -1120
rect 350 -1160 365 -1070
rect 325 -1170 365 -1160
rect 325 -1190 335 -1170
rect 355 -1190 365 -1170
rect 325 -1200 365 -1190
rect 325 -1250 365 -1240
rect 325 -1265 335 -1250
rect 195 -1280 210 -1265
rect 310 -1270 335 -1265
rect 355 -1270 365 -1250
rect 310 -1280 365 -1270
rect 155 -1315 195 -1305
rect 155 -1335 165 -1315
rect 185 -1330 195 -1315
rect 185 -1335 210 -1330
rect 155 -1345 210 -1335
rect 310 -1345 325 -1330
rect 435 -1425 450 -925
rect 550 -955 565 -705
rect 590 -755 630 -745
rect 590 -775 600 -755
rect 620 -775 630 -755
rect 590 -785 630 -775
rect 590 -890 605 -785
rect 760 -810 775 -680
rect 630 -825 645 -810
rect 745 -825 775 -810
rect 590 -900 630 -890
rect 590 -920 600 -900
rect 620 -920 630 -900
rect 590 -930 630 -920
rect 760 -955 775 -825
rect 550 -970 605 -955
rect 630 -970 645 -955
rect 745 -970 775 -955
rect 590 -1325 605 -970
rect 800 -1035 815 -560
rect 760 -1045 815 -1035
rect 760 -1065 770 -1045
rect 790 -1050 815 -1045
rect 790 -1065 800 -1050
rect 760 -1075 800 -1065
rect 630 -1115 645 -1100
rect 745 -1115 840 -1100
rect 760 -1150 800 -1140
rect 760 -1165 770 -1150
rect 630 -1180 645 -1165
rect 745 -1170 770 -1165
rect 790 -1170 800 -1150
rect 745 -1180 800 -1170
rect 825 -1245 840 -1115
rect 650 -1255 840 -1245
rect 650 -1275 660 -1255
rect 680 -1260 840 -1255
rect 680 -1275 690 -1260
rect 650 -1285 690 -1275
rect 590 -1335 630 -1325
rect 590 -1355 600 -1335
rect 620 -1350 630 -1335
rect 620 -1355 645 -1350
rect 590 -1365 645 -1355
rect 745 -1365 760 -1350
rect 760 -1400 800 -1390
rect 760 -1415 770 -1400
rect 410 -1435 450 -1425
rect 630 -1430 645 -1415
rect 745 -1420 770 -1415
rect 790 -1420 800 -1400
rect 745 -1430 800 -1420
rect 410 -1455 420 -1435
rect 440 -1455 450 -1435
rect 410 -1465 450 -1455
<< polycont >>
rect 600 480 620 500
rect 125 300 145 320
rect 335 340 355 360
rect 770 415 790 435
rect 770 335 790 355
rect 335 190 355 210
rect 335 125 355 145
rect 115 -125 135 -105
rect 560 270 580 290
rect 600 165 620 185
rect 600 65 620 85
rect 560 -15 580 5
rect 155 -260 175 -240
rect 115 -385 135 -365
rect 340 -260 360 -240
rect 155 -475 175 -455
rect 400 -360 420 -340
rect 335 -575 355 -555
rect 600 -80 620 -60
rect 810 -35 830 -15
rect 810 -205 830 -185
rect 685 -370 705 -350
rect 750 -410 770 -390
rect 810 -515 830 -495
rect 600 -630 620 -610
rect 560 -695 580 -675
rect 165 -1125 185 -1105
rect 335 -1190 355 -1170
rect 335 -1270 355 -1250
rect 165 -1335 185 -1315
rect 600 -775 620 -755
rect 600 -920 620 -900
rect 770 -1065 790 -1045
rect 770 -1170 790 -1150
rect 660 -1275 680 -1255
rect 600 -1355 620 -1335
rect 770 -1420 790 -1400
rect 420 -1455 440 -1435
<< locali >>
rect 650 545 740 555
rect 650 525 660 545
rect 730 540 740 545
rect 730 525 780 540
rect 650 520 780 525
rect 650 515 740 520
rect 590 500 630 510
rect 590 480 600 500
rect 620 480 630 500
rect 590 470 630 480
rect 215 405 305 415
rect 215 395 225 405
rect 135 385 225 395
rect 295 385 305 405
rect 135 375 305 385
rect 385 410 425 420
rect 135 330 155 375
rect 325 360 365 370
rect 215 340 305 350
rect 215 330 225 340
rect 115 320 155 330
rect 115 300 125 320
rect 145 300 155 320
rect 115 290 155 300
rect 175 320 225 330
rect 295 320 305 340
rect 325 340 335 360
rect 355 340 365 360
rect 325 330 365 340
rect 385 340 395 410
rect 415 340 425 410
rect 385 330 425 340
rect 175 310 305 320
rect 120 -95 140 290
rect 175 -10 195 310
rect 215 275 305 285
rect 215 255 225 275
rect 295 265 305 275
rect 330 265 350 330
rect 550 320 590 410
rect 610 405 630 470
rect 650 480 740 490
rect 650 460 660 480
rect 730 460 740 480
rect 650 450 740 460
rect 760 445 780 520
rect 760 435 800 445
rect 650 415 740 425
rect 650 405 660 415
rect 610 395 660 405
rect 730 395 740 415
rect 760 415 770 435
rect 790 425 800 435
rect 790 415 840 425
rect 760 405 840 415
rect 610 385 740 395
rect 550 290 590 300
rect 550 270 560 290
rect 580 270 590 290
rect 295 255 405 265
rect 215 245 405 255
rect 325 210 365 220
rect 325 200 335 210
rect 215 190 335 200
rect 355 190 365 210
rect 215 170 225 190
rect 295 180 365 190
rect 295 170 305 180
rect 215 160 305 170
rect 325 145 365 155
rect 215 125 305 135
rect 215 105 225 125
rect 295 105 305 125
rect 325 125 335 145
rect 355 125 365 145
rect 325 115 365 125
rect 215 95 305 105
rect 215 60 305 70
rect 215 40 225 60
rect 295 50 305 60
rect 330 50 350 115
rect 385 95 405 245
rect 295 40 350 50
rect 215 30 350 40
rect 175 -20 245 -10
rect 175 -30 215 -20
rect 205 -90 215 -30
rect 235 -90 245 -20
rect 105 -105 145 -95
rect 205 -100 245 -90
rect 270 -20 310 -10
rect 270 -90 280 -20
rect 300 -90 310 -20
rect 270 -100 310 -90
rect 105 -125 115 -105
rect 135 -125 145 -105
rect 105 -135 145 -125
rect 205 -150 245 -140
rect 205 -155 215 -150
rect 85 -175 215 -155
rect 205 -220 215 -175
rect 235 -220 245 -150
rect 205 -230 245 -220
rect 270 -150 310 -140
rect 270 -220 280 -150
rect 300 -220 310 -150
rect 270 -230 310 -220
rect 330 -230 350 30
rect 370 75 405 95
rect 550 260 590 270
rect 550 135 570 260
rect 610 195 630 385
rect 760 355 800 365
rect 760 345 770 355
rect 650 335 770 345
rect 790 335 800 355
rect 650 315 660 335
rect 730 325 800 335
rect 730 315 740 325
rect 650 305 740 315
rect 650 270 740 280
rect 650 250 660 270
rect 730 260 740 270
rect 730 250 780 260
rect 650 240 780 250
rect 590 185 630 195
rect 590 165 600 185
rect 620 165 630 185
rect 590 155 630 165
rect 650 205 740 215
rect 650 185 660 205
rect 730 185 740 205
rect 650 175 740 185
rect 650 135 670 175
rect 550 115 670 135
rect 370 -150 390 75
rect 550 15 570 115
rect 590 85 630 95
rect 590 65 600 85
rect 620 65 630 85
rect 760 75 780 240
rect 590 55 630 65
rect 550 5 590 15
rect 550 -15 560 5
rect 580 -15 590 5
rect 550 -25 590 -15
rect 610 -50 630 55
rect 650 65 780 75
rect 650 45 660 65
rect 730 55 780 65
rect 730 45 740 55
rect 650 35 740 45
rect 820 35 840 405
rect 760 15 840 35
rect 650 0 740 10
rect 650 -20 660 0
rect 730 -20 740 0
rect 650 -30 740 -20
rect 590 -60 630 -50
rect 590 -80 600 -60
rect 620 -70 630 -60
rect 620 -80 740 -70
rect 590 -90 660 -80
rect 650 -100 660 -90
rect 730 -100 740 -80
rect 650 -110 740 -100
rect 650 -145 740 -135
rect 370 -155 450 -150
rect 650 -155 660 -145
rect 370 -170 470 -155
rect 370 -190 390 -170
rect 430 -175 470 -170
rect 540 -165 660 -155
rect 730 -165 740 -145
rect 540 -175 740 -165
rect 370 -210 410 -190
rect 145 -240 185 -230
rect 145 -260 155 -240
rect 175 -250 185 -240
rect 270 -250 290 -230
rect 330 -240 370 -230
rect 330 -250 340 -240
rect 175 -260 290 -250
rect 145 -270 290 -260
rect 310 -260 340 -250
rect 360 -260 370 -240
rect 310 -270 370 -260
rect 310 -290 330 -270
rect 390 -290 410 -210
rect 760 -215 780 15
rect 800 -15 840 -5
rect 800 -35 810 -15
rect 830 -35 840 -15
rect 800 -45 840 -35
rect 820 -155 840 -45
rect 820 -175 850 -155
rect 800 -185 840 -175
rect 800 -205 810 -185
rect 830 -205 840 -185
rect 800 -215 840 -205
rect 650 -225 780 -215
rect 650 -245 660 -225
rect 730 -235 780 -225
rect 730 -245 740 -235
rect 650 -255 740 -245
rect 205 -300 245 -290
rect 205 -315 215 -300
rect 85 -335 215 -315
rect 105 -365 145 -355
rect 105 -385 115 -365
rect 135 -385 145 -365
rect 205 -370 215 -335
rect 235 -370 245 -300
rect 205 -380 245 -370
rect 270 -300 330 -290
rect 270 -370 280 -300
rect 300 -310 330 -300
rect 350 -310 410 -290
rect 650 -290 740 -280
rect 650 -300 660 -290
rect 540 -310 660 -300
rect 730 -310 740 -290
rect 300 -370 310 -310
rect 270 -380 310 -370
rect 105 -395 145 -385
rect 105 -500 125 -395
rect 350 -445 370 -310
rect 430 -330 470 -315
rect 540 -320 740 -310
rect 390 -335 470 -330
rect 390 -340 450 -335
rect 390 -360 400 -340
rect 420 -350 450 -340
rect 675 -350 715 -340
rect 420 -360 430 -350
rect 390 -370 430 -360
rect 675 -370 685 -350
rect 705 -370 715 -350
rect 675 -380 715 -370
rect 760 -380 780 -235
rect 740 -390 780 -380
rect 740 -410 750 -390
rect 770 -410 780 -390
rect 740 -420 780 -410
rect 800 -320 850 -300
rect 800 -445 820 -320
rect 145 -455 245 -445
rect 145 -475 155 -455
rect 175 -465 215 -455
rect 175 -475 185 -465
rect 145 -485 185 -475
rect 105 -520 135 -500
rect 115 -665 135 -520
rect 205 -525 215 -465
rect 235 -525 245 -455
rect 205 -535 245 -525
rect 270 -455 390 -445
rect 270 -525 280 -455
rect 300 -465 390 -455
rect 300 -525 310 -465
rect 370 -505 390 -465
rect 370 -525 405 -505
rect 270 -535 310 -525
rect 325 -555 365 -545
rect 325 -575 335 -555
rect 355 -575 365 -555
rect 325 -585 365 -575
rect 205 -605 245 -595
rect 205 -665 215 -605
rect 115 -675 215 -665
rect 235 -675 245 -605
rect 115 -685 245 -675
rect 270 -605 310 -595
rect 330 -605 350 -585
rect 270 -675 280 -605
rect 300 -625 350 -605
rect 300 -675 310 -625
rect 270 -685 310 -675
rect 330 -670 350 -625
rect 385 -630 405 -525
rect 630 -540 670 -450
rect 740 -465 820 -445
rect 740 -560 760 -465
rect 800 -495 840 -485
rect 800 -515 810 -495
rect 830 -515 840 -495
rect 800 -525 840 -515
rect 550 -580 760 -560
rect 385 -650 435 -630
rect 115 -1305 135 -685
rect 330 -690 395 -670
rect 190 -745 310 -735
rect 190 -765 200 -745
rect 300 -765 310 -745
rect 190 -775 310 -765
rect 190 -810 310 -800
rect 190 -830 200 -810
rect 300 -820 310 -810
rect 300 -830 350 -820
rect 190 -840 350 -830
rect 245 -890 285 -880
rect 245 -960 255 -890
rect 275 -960 285 -890
rect 245 -970 285 -960
rect 215 -1020 305 -1010
rect 215 -1030 225 -1020
rect 175 -1040 225 -1030
rect 295 -1040 305 -1020
rect 175 -1050 305 -1040
rect 175 -1095 195 -1050
rect 330 -1075 350 -840
rect 155 -1105 195 -1095
rect 155 -1125 165 -1105
rect 185 -1125 195 -1105
rect 215 -1085 350 -1075
rect 215 -1105 225 -1085
rect 295 -1095 350 -1085
rect 295 -1105 305 -1095
rect 215 -1115 305 -1105
rect 155 -1135 195 -1125
rect 215 -1150 305 -1140
rect 215 -1170 225 -1150
rect 295 -1160 305 -1150
rect 375 -1160 395 -690
rect 295 -1170 395 -1160
rect 215 -1180 335 -1170
rect 325 -1190 335 -1180
rect 355 -1180 395 -1170
rect 355 -1190 365 -1180
rect 325 -1200 365 -1190
rect 215 -1230 305 -1220
rect 215 -1240 225 -1230
rect 165 -1250 225 -1240
rect 295 -1250 305 -1230
rect 415 -1240 435 -650
rect 550 -665 570 -580
rect 590 -610 630 -600
rect 590 -630 600 -610
rect 620 -620 630 -610
rect 620 -630 740 -620
rect 590 -640 660 -630
rect 550 -675 590 -665
rect 550 -695 560 -675
rect 580 -695 590 -675
rect 550 -705 590 -695
rect 550 -850 570 -705
rect 610 -745 630 -640
rect 650 -650 660 -640
rect 730 -650 740 -630
rect 650 -660 740 -650
rect 650 -695 740 -685
rect 650 -715 660 -695
rect 730 -705 740 -695
rect 820 -705 840 -525
rect 730 -715 840 -705
rect 650 -725 840 -715
rect 590 -755 630 -745
rect 590 -775 600 -755
rect 620 -775 630 -755
rect 590 -785 630 -775
rect 650 -775 780 -765
rect 650 -795 660 -775
rect 730 -785 780 -775
rect 730 -795 740 -785
rect 650 -805 740 -795
rect 650 -840 740 -830
rect 650 -850 660 -840
rect 550 -860 660 -850
rect 730 -860 740 -840
rect 550 -870 740 -860
rect 590 -900 630 -890
rect 590 -920 600 -900
rect 620 -920 630 -900
rect 590 -930 630 -920
rect 610 -955 630 -930
rect 650 -920 740 -910
rect 650 -940 660 -920
rect 730 -940 740 -920
rect 650 -950 740 -940
rect 165 -1260 305 -1250
rect 325 -1250 435 -1240
rect 165 -1305 185 -1260
rect 325 -1270 335 -1250
rect 355 -1260 435 -1250
rect 570 -975 630 -955
rect 570 -1245 590 -975
rect 650 -985 740 -975
rect 650 -995 660 -985
rect 610 -1005 660 -995
rect 730 -1005 740 -985
rect 610 -1015 740 -1005
rect 610 -1120 630 -1015
rect 760 -1035 780 -785
rect 760 -1045 800 -1035
rect 760 -1055 770 -1045
rect 650 -1065 770 -1055
rect 790 -1065 800 -1045
rect 650 -1085 660 -1065
rect 730 -1075 800 -1065
rect 730 -1085 740 -1075
rect 650 -1095 740 -1085
rect 610 -1130 740 -1120
rect 610 -1140 660 -1130
rect 650 -1150 660 -1140
rect 730 -1150 740 -1130
rect 650 -1160 740 -1150
rect 760 -1140 780 -1075
rect 760 -1150 800 -1140
rect 760 -1170 770 -1150
rect 790 -1170 800 -1150
rect 760 -1180 800 -1170
rect 650 -1195 740 -1185
rect 650 -1215 660 -1195
rect 730 -1215 740 -1195
rect 820 -1200 840 -725
rect 650 -1225 740 -1215
rect 760 -1220 840 -1200
rect 650 -1245 670 -1225
rect 570 -1255 690 -1245
rect 355 -1270 365 -1260
rect 570 -1265 660 -1255
rect 325 -1280 365 -1270
rect 650 -1275 660 -1265
rect 680 -1275 690 -1255
rect 215 -1295 305 -1285
rect 115 -1315 195 -1305
rect 115 -1325 165 -1315
rect 155 -1335 165 -1325
rect 185 -1335 195 -1315
rect 215 -1315 225 -1295
rect 295 -1315 305 -1295
rect 215 -1325 305 -1315
rect 155 -1345 195 -1335
rect 330 -1350 350 -1280
rect 650 -1285 690 -1275
rect 650 -1315 740 -1305
rect 215 -1360 350 -1350
rect 215 -1380 225 -1360
rect 295 -1370 350 -1360
rect 590 -1335 630 -1325
rect 590 -1355 600 -1335
rect 620 -1355 630 -1335
rect 650 -1335 660 -1315
rect 730 -1325 740 -1315
rect 760 -1325 780 -1220
rect 730 -1335 780 -1325
rect 650 -1345 780 -1335
rect 590 -1365 630 -1355
rect 295 -1380 305 -1370
rect 215 -1390 305 -1380
rect 410 -1435 450 -1425
rect 410 -1455 420 -1435
rect 440 -1455 450 -1435
rect 610 -1435 630 -1365
rect 650 -1380 740 -1370
rect 650 -1400 660 -1380
rect 730 -1400 740 -1380
rect 650 -1410 740 -1400
rect 760 -1390 780 -1345
rect 760 -1400 800 -1390
rect 760 -1420 770 -1400
rect 790 -1420 800 -1400
rect 760 -1430 800 -1420
rect 610 -1445 740 -1435
rect 610 -1455 660 -1445
rect 410 -1465 450 -1455
rect 650 -1465 660 -1455
rect 730 -1465 740 -1445
rect 650 -1475 740 -1465
<< viali >>
rect 395 340 415 410
rect 225 105 295 125
rect 280 -90 300 -20
rect 200 -765 300 -745
rect 255 -960 275 -890
rect 225 -1315 295 -1295
rect 420 -1455 440 -1435
<< metal1 >>
rect 85 410 470 425
rect 85 340 395 410
rect 415 340 470 410
rect 85 125 470 340
rect 85 105 225 125
rect 295 105 470 125
rect 85 -20 470 105
rect 85 -90 280 -20
rect 300 -90 470 -20
rect 85 -105 470 -90
rect 85 -745 470 -730
rect 85 -765 200 -745
rect 300 -765 470 -745
rect 85 -890 470 -765
rect 85 -960 255 -890
rect 275 -960 470 -890
rect 85 -1295 470 -960
rect 85 -1315 225 -1295
rect 295 -1315 470 -1295
rect 85 -1395 470 -1315
rect 85 -1435 470 -1425
rect 85 -1455 420 -1435
rect 440 -1455 470 -1435
rect 85 -1465 470 -1455
<< labels >>
rlabel locali 85 -165 85 -165 7 D
rlabel locali 85 -325 85 -325 7 D_BAR
rlabel locali 470 -165 470 -165 3 Q
rlabel locali 470 -325 470 -325 3 Q_BAR
rlabel metal1 85 155 85 155 7 VP
rlabel metal1 85 -1270 85 -1270 7 VN
rlabel metal1 85 -1445 85 -1445 7 CLK
<< end >>
