magic
tech sky130A
timestamp 1695522088
<< nwell >>
rect -70 -145 400 340
<< nmos >>
rect 0 -410 15 -310
rect 65 -410 80 -310
rect 250 -410 265 -310
rect 250 -545 265 -445
rect -15 -645 120 -630
rect -15 -710 120 -695
rect 250 -755 265 -655
rect 315 -755 330 -655
rect -15 -775 120 -760
<< pmos >>
rect 0 220 15 320
rect 65 220 80 320
rect 195 215 295 230
rect 0 10 15 110
rect 0 -125 15 -25
rect 250 -125 265 -25
rect 315 -125 330 -25
<< ndiff >>
rect -50 -325 0 -310
rect -50 -395 -35 -325
rect -15 -395 0 -325
rect -50 -410 0 -395
rect 15 -325 65 -310
rect 15 -395 30 -325
rect 50 -395 65 -325
rect 15 -410 65 -395
rect 80 -325 130 -310
rect 80 -395 95 -325
rect 115 -395 130 -325
rect 80 -410 130 -395
rect 200 -325 250 -310
rect 200 -395 215 -325
rect 235 -395 250 -325
rect 200 -410 250 -395
rect 265 -325 315 -310
rect 265 -395 280 -325
rect 300 -395 315 -325
rect 265 -410 315 -395
rect 200 -460 250 -445
rect 200 -530 215 -460
rect 235 -530 250 -460
rect 200 -545 250 -530
rect 265 -460 315 -445
rect 265 -530 280 -460
rect 300 -530 315 -460
rect 265 -545 315 -530
rect -15 -595 120 -580
rect -15 -615 0 -595
rect 105 -615 120 -595
rect -15 -630 120 -615
rect -15 -660 120 -645
rect -15 -680 0 -660
rect 105 -680 120 -660
rect -15 -695 120 -680
rect -15 -725 120 -710
rect -15 -745 0 -725
rect 105 -745 120 -725
rect -15 -760 120 -745
rect 200 -670 250 -655
rect 200 -740 215 -670
rect 235 -740 250 -670
rect 200 -755 250 -740
rect 265 -670 315 -655
rect 265 -740 280 -670
rect 300 -740 315 -670
rect 265 -755 315 -740
rect 330 -670 380 -655
rect 330 -740 345 -670
rect 365 -740 380 -670
rect 330 -755 380 -740
rect -15 -790 120 -775
rect -15 -810 0 -790
rect 105 -810 120 -790
rect -15 -825 120 -810
<< pdiff >>
rect -50 305 0 320
rect -50 235 -35 305
rect -15 235 0 305
rect -50 220 0 235
rect 15 305 65 320
rect 15 235 30 305
rect 50 235 65 305
rect 15 220 65 235
rect 80 305 130 320
rect 80 235 95 305
rect 115 235 130 305
rect 80 220 130 235
rect 195 265 295 280
rect 195 245 210 265
rect 280 245 295 265
rect 195 230 295 245
rect -50 95 0 110
rect -50 25 -35 95
rect -15 25 0 95
rect -50 10 0 25
rect 15 95 65 110
rect 15 25 30 95
rect 50 25 65 95
rect 15 10 65 25
rect -50 -40 0 -25
rect -50 -110 -35 -40
rect -15 -110 0 -40
rect -50 -125 0 -110
rect 15 -40 65 -25
rect 15 -110 30 -40
rect 50 -110 65 -40
rect 15 -125 65 -110
rect 195 200 295 215
rect 195 180 210 200
rect 280 180 295 200
rect 195 165 295 180
rect 200 -40 250 -25
rect 200 -110 215 -40
rect 235 -110 250 -40
rect 200 -125 250 -110
rect 265 -40 315 -25
rect 265 -110 280 -40
rect 300 -110 315 -40
rect 265 -125 315 -110
rect 330 -40 380 -25
rect 330 -110 345 -40
rect 365 -110 380 -40
rect 330 -125 380 -110
<< ndiffc >>
rect -35 -395 -15 -325
rect 30 -395 50 -325
rect 95 -395 115 -325
rect 215 -395 235 -325
rect 280 -395 300 -325
rect 215 -530 235 -460
rect 280 -530 300 -460
rect 0 -615 105 -595
rect 0 -680 105 -660
rect 0 -745 105 -725
rect 215 -740 235 -670
rect 280 -740 300 -670
rect 345 -740 365 -670
rect 0 -810 105 -790
<< pdiffc >>
rect -35 235 -15 305
rect 30 235 50 305
rect 95 235 115 305
rect 210 245 280 265
rect -35 25 -15 95
rect 30 25 50 95
rect -35 -110 -15 -40
rect 30 -110 50 -40
rect 210 180 280 200
rect 215 -110 235 -40
rect 280 -110 300 -40
rect 345 -110 365 -40
<< psubdiff >>
rect 70 -515 170 -500
rect 70 -535 85 -515
rect 155 -535 170 -515
rect 70 -550 170 -535
<< nsubdiff >>
rect 245 120 345 135
rect 245 100 260 120
rect 330 100 345 120
rect 245 85 345 100
<< psubdiffcont >>
rect 85 -535 155 -515
<< nsubdiffcont >>
rect 260 100 330 120
<< poly >>
rect 0 365 40 375
rect 0 345 10 365
rect 30 345 40 365
rect 0 335 40 345
rect 0 320 15 335
rect 65 320 80 335
rect 0 205 15 220
rect 65 205 80 220
rect 165 215 195 230
rect 295 215 310 230
rect 65 195 105 205
rect 65 175 75 195
rect 95 175 105 195
rect 65 165 105 175
rect 0 110 15 125
rect 0 -25 15 10
rect 0 -190 15 -125
rect 165 -190 180 215
rect 250 60 290 70
rect 250 40 260 60
rect 280 40 290 60
rect 250 30 290 40
rect 395 45 435 55
rect 250 -25 265 30
rect 395 25 405 45
rect 425 25 435 45
rect 395 15 435 25
rect 315 -25 330 -10
rect 250 -140 265 -125
rect 315 -140 330 -125
rect 395 -135 410 15
rect 295 -155 330 -140
rect 375 -150 410 -135
rect 295 -165 310 -155
rect 270 -175 310 -165
rect -50 -205 245 -190
rect 270 -195 280 -175
rect 300 -195 310 -175
rect 270 -205 310 -195
rect 150 -240 190 -230
rect 150 -255 160 -240
rect 40 -260 160 -255
rect 180 -260 190 -240
rect 230 -235 245 -205
rect 310 -235 350 -230
rect 230 -240 350 -235
rect 230 -250 320 -240
rect 40 -265 190 -260
rect 40 -285 50 -265
rect 70 -270 190 -265
rect 70 -285 80 -270
rect 40 -295 80 -285
rect 0 -310 15 -295
rect 65 -310 80 -295
rect 250 -310 265 -250
rect 310 -260 320 -250
rect 340 -260 350 -240
rect 310 -270 350 -260
rect 375 -295 390 -150
rect 435 -205 455 -190
rect 435 -230 450 -205
rect 415 -240 455 -230
rect 415 -260 425 -240
rect 445 -260 455 -240
rect 415 -270 455 -260
rect 330 -310 390 -295
rect 0 -465 15 -410
rect 65 -425 80 -410
rect 250 -445 265 -410
rect 0 -475 40 -465
rect 0 -495 10 -475
rect 30 -495 40 -475
rect 0 -505 40 -495
rect 250 -580 265 -545
rect 130 -595 265 -580
rect 130 -630 145 -595
rect 330 -600 345 -310
rect -30 -645 -15 -630
rect 120 -645 145 -630
rect 290 -610 345 -600
rect 290 -630 300 -610
rect 320 -615 345 -610
rect 320 -630 330 -615
rect 290 -640 330 -630
rect 130 -695 145 -645
rect 250 -655 265 -640
rect 315 -655 330 -640
rect -30 -710 -15 -695
rect 120 -710 145 -695
rect 130 -760 145 -710
rect -30 -775 -15 -760
rect 120 -775 145 -760
rect 250 -770 265 -755
rect 315 -770 330 -755
rect 250 -780 290 -770
rect 250 -800 260 -780
rect 280 -800 290 -780
rect 250 -810 290 -800
<< polycont >>
rect 10 345 30 365
rect 75 175 95 195
rect 260 40 280 60
rect 405 25 425 45
rect 280 -195 300 -175
rect 160 -260 180 -240
rect 50 -285 70 -265
rect 320 -260 340 -240
rect 425 -260 445 -240
rect 10 -495 30 -475
rect 300 -630 320 -610
rect 260 -800 280 -780
<< locali >>
rect 0 365 40 375
rect 0 345 10 365
rect 30 355 40 365
rect 30 345 125 355
rect 0 335 125 345
rect 105 315 125 335
rect -45 305 -5 315
rect -45 235 -35 305
rect -15 235 -5 305
rect -45 225 -5 235
rect 20 305 60 315
rect 20 235 30 305
rect 50 235 60 305
rect 20 225 60 235
rect 85 305 125 315
rect 85 235 95 305
rect 115 245 125 305
rect 200 265 290 275
rect 200 245 210 265
rect 280 245 290 265
rect 115 235 150 245
rect 200 235 290 245
rect 85 225 150 235
rect -25 205 -5 225
rect -25 195 105 205
rect -25 185 75 195
rect 25 105 45 185
rect 65 175 75 185
rect 95 175 105 195
rect 65 165 105 175
rect -45 95 -5 105
rect -45 35 -35 95
rect -50 25 -35 35
rect -15 25 -5 95
rect -50 15 -5 25
rect 20 95 60 105
rect 20 25 30 95
rect 50 25 60 95
rect 20 15 60 25
rect -45 -40 -5 -30
rect -45 -100 -35 -40
rect -50 -110 -35 -100
rect -15 -110 -5 -40
rect -50 -120 -5 -110
rect 20 -40 60 -30
rect 20 -110 30 -40
rect 50 -110 60 -40
rect 20 -120 60 -110
rect 40 -255 60 -120
rect 85 -215 105 165
rect 130 -150 150 225
rect 200 200 290 210
rect 200 180 210 200
rect 280 180 290 200
rect 200 170 290 180
rect 200 10 220 170
rect 250 120 340 130
rect 250 100 260 120
rect 330 100 340 120
rect 250 90 340 100
rect 250 60 290 70
rect 250 40 260 60
rect 280 50 290 60
rect 395 50 435 55
rect 280 45 435 50
rect 280 40 405 45
rect 250 30 405 40
rect 200 -10 290 10
rect 270 -30 290 -10
rect 355 -30 375 30
rect 395 25 405 30
rect 425 35 435 45
rect 425 25 455 35
rect 395 15 455 25
rect 205 -40 245 -30
rect 205 -110 215 -40
rect 235 -110 245 -40
rect 205 -120 245 -110
rect 270 -40 310 -30
rect 270 -110 280 -40
rect 300 -110 310 -40
rect 270 -120 310 -110
rect 335 -40 375 -30
rect 335 -110 345 -40
rect 365 -110 375 -40
rect 335 -120 375 -110
rect 405 -120 455 -100
rect 225 -140 245 -120
rect 130 -170 170 -150
rect 225 -160 290 -140
rect 85 -235 125 -215
rect 40 -265 80 -255
rect 40 -275 50 -265
rect -25 -285 50 -275
rect 70 -285 80 -265
rect -25 -295 80 -285
rect -25 -315 -5 -295
rect 105 -315 125 -235
rect 150 -230 170 -170
rect 270 -165 290 -160
rect 405 -165 425 -120
rect 270 -175 425 -165
rect 270 -195 280 -175
rect 300 -185 425 -175
rect 300 -195 310 -185
rect 270 -205 310 -195
rect 150 -240 190 -230
rect 150 -260 160 -240
rect 180 -250 190 -240
rect 180 -260 225 -250
rect 150 -270 225 -260
rect -45 -325 -5 -315
rect -45 -395 -35 -325
rect -15 -395 -5 -325
rect -45 -405 -5 -395
rect 20 -325 60 -315
rect 20 -395 30 -325
rect 50 -395 60 -325
rect 20 -405 60 -395
rect 85 -325 125 -315
rect 85 -395 95 -325
rect 115 -395 125 -325
rect 85 -405 125 -395
rect 205 -315 225 -270
rect 270 -315 290 -205
rect 310 -240 455 -230
rect 310 -260 320 -240
rect 340 -250 425 -240
rect 340 -260 350 -250
rect 310 -270 350 -260
rect 415 -260 425 -250
rect 445 -260 455 -240
rect 415 -270 455 -260
rect 205 -325 245 -315
rect 205 -395 215 -325
rect 235 -395 245 -325
rect 205 -405 245 -395
rect 270 -325 310 -315
rect 270 -395 280 -325
rect 300 -385 310 -325
rect 300 -395 375 -385
rect 270 -405 375 -395
rect 20 -425 40 -405
rect -50 -445 40 -425
rect -50 -585 -30 -445
rect 105 -465 125 -405
rect 205 -460 245 -450
rect 205 -465 215 -460
rect 0 -475 215 -465
rect 0 -495 10 -475
rect 30 -485 215 -475
rect 30 -495 40 -485
rect 0 -505 40 -495
rect 75 -515 165 -505
rect 75 -535 85 -515
rect 155 -535 165 -515
rect 75 -545 165 -535
rect 205 -530 215 -485
rect 235 -530 245 -460
rect 205 -540 245 -530
rect 270 -460 310 -450
rect 270 -530 280 -460
rect 300 -530 310 -460
rect 270 -540 310 -530
rect -50 -595 115 -585
rect -50 -605 0 -595
rect -50 -715 -30 -605
rect -10 -615 0 -605
rect 105 -615 115 -595
rect -10 -625 115 -615
rect 290 -600 310 -540
rect 290 -610 330 -600
rect 290 -620 300 -610
rect 225 -630 300 -620
rect 320 -630 330 -610
rect 225 -640 330 -630
rect -10 -660 115 -650
rect 225 -660 245 -640
rect 355 -660 375 -405
rect -10 -680 0 -660
rect 105 -680 115 -660
rect -10 -690 115 -680
rect 205 -670 245 -660
rect -50 -725 115 -715
rect -50 -735 0 -725
rect -10 -745 0 -735
rect 105 -745 115 -725
rect -10 -755 115 -745
rect 205 -740 215 -670
rect 235 -740 245 -670
rect 205 -750 245 -740
rect 270 -670 310 -660
rect 270 -740 280 -670
rect 300 -740 310 -670
rect 270 -750 310 -740
rect 335 -670 375 -660
rect 335 -740 345 -670
rect 365 -740 375 -670
rect 335 -750 375 -740
rect 355 -770 375 -750
rect 250 -780 375 -770
rect -10 -790 115 -780
rect -10 -810 0 -790
rect 105 -810 115 -790
rect 250 -800 260 -780
rect 280 -790 375 -780
rect 280 -800 290 -790
rect 250 -810 290 -800
rect -10 -820 115 -810
<< end >>
