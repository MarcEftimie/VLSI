magic
tech sky130A
timestamp 1695595790
<< nmos >>
rect 210 325 310 340
rect 210 260 310 275
rect 210 115 310 130
rect 210 50 310 65
rect 250 -130 265 -30
rect 250 -260 265 -160
rect 250 -410 265 -310
rect 250 -540 265 -440
rect 250 -690 265 -590
rect 185 -795 315 -780
rect 185 -860 315 -845
rect 185 -925 315 -910
rect 210 -1070 310 -1055
rect 210 -1135 310 -1120
rect 210 -1280 310 -1265
rect 210 -1345 310 -1330
<< ndiff >>
rect 210 375 310 390
rect 210 355 225 375
rect 295 355 310 375
rect 210 340 310 355
rect 210 310 310 325
rect 210 290 225 310
rect 295 290 310 310
rect 210 275 310 290
rect 210 245 310 260
rect 210 225 225 245
rect 295 225 310 245
rect 210 210 310 225
rect 210 165 310 180
rect 210 145 225 165
rect 295 145 310 165
rect 210 130 310 145
rect 210 100 310 115
rect 210 80 225 100
rect 295 80 310 100
rect 210 65 310 80
rect 210 35 310 50
rect 210 15 225 35
rect 295 15 310 35
rect 210 0 310 15
rect 200 -45 250 -30
rect 200 -115 215 -45
rect 235 -115 250 -45
rect 200 -130 250 -115
rect 265 -45 315 -30
rect 265 -115 280 -45
rect 300 -115 315 -45
rect 265 -130 315 -115
rect 200 -175 250 -160
rect 200 -245 215 -175
rect 235 -245 250 -175
rect 200 -260 250 -245
rect 265 -175 315 -160
rect 265 -245 280 -175
rect 300 -245 315 -175
rect 265 -260 315 -245
rect 200 -325 250 -310
rect 200 -395 215 -325
rect 235 -395 250 -325
rect 200 -410 250 -395
rect 265 -325 315 -310
rect 265 -395 280 -325
rect 300 -395 315 -325
rect 265 -410 315 -395
rect 200 -455 250 -440
rect 200 -525 215 -455
rect 235 -525 250 -455
rect 200 -540 250 -525
rect 265 -455 315 -440
rect 265 -525 280 -455
rect 300 -525 315 -455
rect 265 -540 315 -525
rect 200 -605 250 -590
rect 200 -675 215 -605
rect 235 -675 250 -605
rect 200 -690 250 -675
rect 265 -605 315 -590
rect 265 -675 280 -605
rect 300 -675 315 -605
rect 265 -690 315 -675
rect 185 -745 315 -730
rect 185 -765 200 -745
rect 300 -765 315 -745
rect 185 -780 315 -765
rect 185 -810 315 -795
rect 185 -830 200 -810
rect 300 -830 315 -810
rect 185 -845 315 -830
rect 185 -875 315 -860
rect 185 -895 200 -875
rect 300 -895 315 -875
rect 185 -910 315 -895
rect 185 -940 315 -925
rect 185 -960 200 -940
rect 300 -960 315 -940
rect 185 -975 315 -960
rect 210 -1020 310 -1005
rect 210 -1040 225 -1020
rect 295 -1040 310 -1020
rect 210 -1055 310 -1040
rect 210 -1085 310 -1070
rect 210 -1105 225 -1085
rect 295 -1105 310 -1085
rect 210 -1120 310 -1105
rect 210 -1150 310 -1135
rect 210 -1170 225 -1150
rect 295 -1170 310 -1150
rect 210 -1185 310 -1170
rect 210 -1230 310 -1215
rect 210 -1250 225 -1230
rect 295 -1250 310 -1230
rect 210 -1265 310 -1250
rect 210 -1295 310 -1280
rect 210 -1315 225 -1295
rect 295 -1315 310 -1295
rect 210 -1330 310 -1315
rect 210 -1360 310 -1345
rect 210 -1380 225 -1360
rect 295 -1380 310 -1360
rect 210 -1395 310 -1380
<< ndiffc >>
rect 225 355 295 375
rect 225 290 295 310
rect 225 225 295 245
rect 225 145 295 165
rect 225 80 295 100
rect 225 15 295 35
rect 215 -115 235 -45
rect 280 -115 300 -45
rect 215 -245 235 -175
rect 280 -245 300 -175
rect 215 -395 235 -325
rect 280 -395 300 -325
rect 215 -525 235 -455
rect 280 -525 300 -455
rect 215 -675 235 -605
rect 280 -675 300 -605
rect 200 -765 300 -745
rect 200 -830 300 -810
rect 200 -895 300 -875
rect 200 -960 300 -940
rect 225 -1040 295 -1020
rect 225 -1105 295 -1085
rect 225 -1170 295 -1150
rect 225 -1250 295 -1230
rect 225 -1315 295 -1295
rect 225 -1380 295 -1360
<< poly >>
rect 195 325 210 340
rect 310 330 365 340
rect 310 325 335 330
rect 325 310 335 325
rect 355 310 365 330
rect 325 300 365 310
rect 155 265 210 275
rect 155 245 165 265
rect 185 260 210 265
rect 310 260 405 275
rect 185 245 195 260
rect 155 235 195 245
rect 155 185 195 195
rect 155 165 165 185
rect 185 165 195 185
rect 155 155 195 165
rect 155 65 170 155
rect 195 115 210 130
rect 310 120 365 130
rect 310 115 335 120
rect 325 100 335 115
rect 355 100 365 120
rect 325 90 365 100
rect 155 50 210 65
rect 310 50 325 65
rect 105 -130 145 -120
rect 105 -150 115 -130
rect 135 -150 145 -130
rect 105 -160 145 -150
rect 105 -380 120 -160
rect 170 -255 185 50
rect 250 -30 265 -15
rect 250 -160 265 -130
rect 145 -265 185 -255
rect 390 -205 405 260
rect 390 -220 410 -205
rect 145 -285 155 -265
rect 175 -285 185 -265
rect 145 -295 185 -285
rect 105 -390 145 -380
rect 105 -410 115 -390
rect 135 -410 145 -390
rect 105 -420 145 -410
rect 170 -445 185 -295
rect 250 -310 265 -260
rect 330 -265 370 -255
rect 330 -285 340 -265
rect 360 -285 370 -265
rect 330 -295 370 -285
rect 250 -440 265 -410
rect 145 -455 185 -445
rect 145 -475 155 -455
rect 175 -475 185 -455
rect 145 -485 185 -475
rect 170 -700 185 -485
rect 250 -590 265 -540
rect 335 -545 350 -295
rect 395 -305 410 -220
rect 390 -320 410 -305
rect 390 -355 405 -320
rect 390 -365 430 -355
rect 390 -385 400 -365
rect 420 -385 430 -365
rect 390 -395 430 -385
rect 325 -555 365 -545
rect 325 -575 335 -555
rect 355 -575 365 -555
rect 325 -585 365 -575
rect 130 -715 185 -700
rect 250 -705 265 -690
rect 130 -955 145 -715
rect 250 -720 345 -705
rect 330 -780 345 -720
rect 170 -795 185 -780
rect 315 -795 345 -780
rect 330 -845 345 -795
rect 170 -860 185 -845
rect 315 -860 345 -845
rect 330 -910 345 -860
rect 170 -925 185 -910
rect 315 -925 450 -910
rect 130 -970 170 -955
rect 155 -1095 170 -970
rect 370 -1040 410 -1030
rect 370 -1055 380 -1040
rect 195 -1070 210 -1055
rect 310 -1060 380 -1055
rect 400 -1060 410 -1040
rect 310 -1070 410 -1060
rect 155 -1105 195 -1095
rect 155 -1125 165 -1105
rect 185 -1120 195 -1105
rect 185 -1125 210 -1120
rect 155 -1135 210 -1125
rect 310 -1135 325 -1120
rect 325 -1250 365 -1240
rect 325 -1265 335 -1250
rect 195 -1280 210 -1265
rect 310 -1270 335 -1265
rect 355 -1270 365 -1250
rect 310 -1280 365 -1270
rect 155 -1315 195 -1305
rect 155 -1335 165 -1315
rect 185 -1330 195 -1315
rect 185 -1335 210 -1330
rect 155 -1345 210 -1335
rect 310 -1345 325 -1330
rect 435 -1430 450 -925
rect 410 -1440 450 -1430
rect 410 -1460 420 -1440
rect 440 -1460 450 -1440
rect 410 -1470 450 -1460
<< polycont >>
rect 335 310 355 330
rect 165 245 185 265
rect 165 165 185 185
rect 335 100 355 120
rect 115 -150 135 -130
rect 155 -285 175 -265
rect 115 -410 135 -390
rect 340 -285 360 -265
rect 155 -475 175 -455
rect 400 -385 420 -365
rect 335 -575 355 -555
rect 380 -1060 400 -1040
rect 165 -1125 185 -1105
rect 335 -1270 355 -1250
rect 165 -1335 185 -1315
rect 420 -1460 440 -1440
<< locali >>
rect 215 375 305 385
rect 215 365 225 375
rect 165 355 225 365
rect 295 355 305 375
rect 165 345 305 355
rect 165 275 185 345
rect 325 330 365 340
rect 215 310 305 320
rect 215 290 225 310
rect 295 290 305 310
rect 325 310 335 330
rect 355 310 365 330
rect 325 300 365 310
rect 215 280 305 290
rect 155 265 195 275
rect 155 255 165 265
rect 115 245 165 255
rect 185 245 195 265
rect 115 235 195 245
rect 215 245 305 255
rect 115 -120 135 235
rect 215 225 225 245
rect 295 235 305 245
rect 330 235 350 300
rect 295 225 390 235
rect 215 215 390 225
rect 155 185 195 195
rect 155 165 165 185
rect 185 175 195 185
rect 185 165 305 175
rect 155 155 225 165
rect 215 145 225 155
rect 295 145 305 165
rect 370 170 390 215
rect 370 150 405 170
rect 215 135 305 145
rect 325 120 365 130
rect 215 100 305 110
rect 215 90 225 100
rect 175 80 225 90
rect 295 80 305 100
rect 325 100 335 120
rect 355 100 365 120
rect 325 90 365 100
rect 175 70 305 80
rect 175 -35 195 70
rect 215 35 305 45
rect 215 15 225 35
rect 295 25 305 35
rect 330 25 350 90
rect 385 70 405 150
rect 295 15 350 25
rect 215 5 350 15
rect 175 -45 245 -35
rect 175 -55 215 -45
rect 205 -115 215 -55
rect 235 -115 245 -45
rect 105 -130 145 -120
rect 205 -125 245 -115
rect 270 -45 310 -35
rect 270 -115 280 -45
rect 300 -115 310 -45
rect 270 -125 310 -115
rect 105 -150 115 -130
rect 135 -150 145 -130
rect 105 -160 145 -150
rect 205 -175 245 -165
rect 205 -180 215 -175
rect 85 -200 215 -180
rect 205 -245 215 -200
rect 235 -245 245 -175
rect 205 -255 245 -245
rect 270 -175 310 -165
rect 270 -245 280 -175
rect 300 -245 310 -175
rect 270 -255 310 -245
rect 330 -255 350 5
rect 370 50 405 70
rect 370 -175 390 50
rect 370 -180 450 -175
rect 370 -195 465 -180
rect 370 -215 390 -195
rect 430 -200 465 -195
rect 370 -235 410 -215
rect 145 -265 185 -255
rect 145 -285 155 -265
rect 175 -275 185 -265
rect 270 -275 290 -255
rect 330 -265 370 -255
rect 330 -275 340 -265
rect 175 -285 290 -275
rect 145 -295 290 -285
rect 310 -285 340 -275
rect 360 -285 370 -265
rect 310 -295 370 -285
rect 310 -315 330 -295
rect 390 -315 410 -235
rect 205 -325 245 -315
rect 205 -340 215 -325
rect 85 -360 215 -340
rect 105 -390 145 -380
rect 105 -410 115 -390
rect 135 -410 145 -390
rect 205 -395 215 -360
rect 235 -395 245 -325
rect 205 -405 245 -395
rect 270 -325 330 -315
rect 270 -395 280 -325
rect 300 -335 330 -325
rect 350 -335 410 -315
rect 300 -395 310 -335
rect 270 -405 310 -395
rect 105 -420 145 -410
rect 105 -500 125 -420
rect 350 -445 370 -335
rect 430 -355 470 -340
rect 390 -360 470 -355
rect 390 -365 450 -360
rect 390 -385 400 -365
rect 420 -375 450 -365
rect 420 -385 430 -375
rect 390 -395 430 -385
rect 145 -455 245 -445
rect 145 -475 155 -455
rect 175 -465 215 -455
rect 175 -475 185 -465
rect 145 -485 185 -475
rect 105 -520 135 -500
rect 115 -665 135 -520
rect 205 -525 215 -465
rect 235 -525 245 -455
rect 205 -535 245 -525
rect 270 -455 390 -445
rect 270 -525 280 -455
rect 300 -465 390 -455
rect 300 -525 310 -465
rect 370 -505 390 -465
rect 370 -525 405 -505
rect 270 -535 310 -525
rect 325 -555 365 -545
rect 325 -575 335 -555
rect 355 -575 365 -555
rect 325 -585 365 -575
rect 205 -605 245 -595
rect 205 -665 215 -605
rect 115 -675 215 -665
rect 235 -675 245 -605
rect 115 -685 245 -675
rect 270 -605 310 -595
rect 330 -605 350 -585
rect 270 -675 280 -605
rect 300 -625 350 -605
rect 300 -675 310 -625
rect 270 -685 310 -675
rect 330 -670 350 -625
rect 385 -630 405 -525
rect 385 -650 435 -630
rect 115 -1155 135 -685
rect 330 -690 395 -670
rect 190 -745 310 -735
rect 190 -765 200 -745
rect 300 -765 310 -745
rect 190 -775 310 -765
rect 190 -810 310 -800
rect 190 -830 200 -810
rect 300 -820 310 -810
rect 300 -830 350 -820
rect 190 -840 350 -830
rect 190 -875 310 -865
rect 190 -895 200 -875
rect 300 -895 310 -875
rect 190 -905 310 -895
rect 330 -930 350 -840
rect 190 -940 350 -930
rect 190 -960 200 -940
rect 300 -950 350 -940
rect 300 -960 310 -950
rect 190 -970 310 -960
rect 215 -1020 305 -1010
rect 215 -1030 225 -1020
rect 165 -1040 225 -1030
rect 295 -1040 305 -1020
rect 165 -1050 305 -1040
rect 165 -1095 185 -1050
rect 330 -1075 350 -950
rect 375 -1030 395 -690
rect 415 -990 435 -650
rect 415 -1010 450 -990
rect 370 -1040 410 -1030
rect 370 -1060 380 -1040
rect 400 -1060 410 -1040
rect 370 -1070 410 -1060
rect 215 -1085 350 -1075
rect 155 -1105 195 -1095
rect 155 -1125 165 -1105
rect 185 -1125 195 -1105
rect 215 -1105 225 -1085
rect 295 -1095 350 -1085
rect 295 -1105 305 -1095
rect 215 -1115 305 -1105
rect 155 -1135 195 -1125
rect 375 -1140 395 -1070
rect 430 -1090 450 -1010
rect 215 -1150 395 -1140
rect 115 -1175 145 -1155
rect 125 -1240 145 -1175
rect 215 -1170 225 -1150
rect 295 -1160 395 -1150
rect 415 -1110 450 -1090
rect 295 -1170 305 -1160
rect 215 -1180 305 -1170
rect 415 -1180 435 -1110
rect 370 -1200 435 -1180
rect 215 -1230 305 -1220
rect 215 -1240 225 -1230
rect 125 -1250 225 -1240
rect 295 -1250 305 -1230
rect 370 -1240 390 -1200
rect 125 -1260 305 -1250
rect 325 -1250 390 -1240
rect 165 -1305 185 -1260
rect 325 -1270 335 -1250
rect 355 -1260 390 -1250
rect 355 -1270 365 -1260
rect 325 -1280 365 -1270
rect 215 -1295 305 -1285
rect 155 -1315 195 -1305
rect 155 -1335 165 -1315
rect 185 -1335 195 -1315
rect 215 -1315 225 -1295
rect 295 -1315 305 -1295
rect 215 -1325 305 -1315
rect 155 -1345 195 -1335
rect 330 -1350 350 -1280
rect 215 -1360 350 -1350
rect 215 -1380 225 -1360
rect 295 -1370 350 -1360
rect 295 -1380 305 -1370
rect 215 -1390 305 -1380
rect 410 -1440 450 -1430
rect 410 -1460 420 -1440
rect 440 -1460 450 -1440
rect 410 -1470 450 -1460
<< end >>
