magic
tech sky130A
timestamp 1697393108
<< nwell >>
rect -7020 1705 -6970 2895
rect -3410 1510 -3200 2895
<< pmos >>
rect -3320 1570 -3270 2770
<< pdiff >>
rect -3370 2755 -3320 2770
rect -3370 1585 -3355 2755
rect -3335 1585 -3320 2755
rect -3370 1570 -3320 1585
rect -3270 2755 -3220 2770
rect -3270 1585 -3255 2755
rect -3235 1585 -3220 2755
rect -3270 1570 -3220 1585
<< pdiffc >>
rect -3355 1585 -3335 2755
rect -3255 1585 -3235 2755
<< poly >>
rect -4720 2940 -4680 2950
rect -4720 2920 -4710 2940
rect -4690 2920 -4680 2940
rect -4720 2910 -4680 2920
rect -4720 2890 -4705 2910
rect -5200 2875 -4705 2890
rect -3320 2815 -3270 2825
rect -3320 2795 -3310 2815
rect -3290 2795 -3270 2815
rect -3320 2770 -3270 2795
rect -3320 1555 -3270 1570
rect -7620 275 -7580 285
rect -7620 255 -7610 275
rect -7590 255 -7580 275
rect -7620 245 -7580 255
rect -7095 275 -7055 285
rect -7095 255 -7085 275
rect -7065 255 -7055 275
rect -7095 245 -7055 255
rect -7620 95 -7605 245
rect -7095 95 -7080 245
rect -6780 145 -6740 155
rect -6655 145 -6615 155
rect -6780 125 -6770 145
rect -6750 130 -6645 145
rect -6750 125 -6740 130
rect -6780 115 -6740 125
rect -6655 125 -6645 130
rect -6625 125 -6615 145
rect -6655 115 -6615 125
rect -7620 85 -7580 95
rect -7620 65 -7610 85
rect -7590 65 -7580 85
rect -7620 55 -7580 65
rect -7095 85 -7055 95
rect -7095 65 -7085 85
rect -7065 65 -7055 85
rect -7095 55 -7055 65
<< polycont >>
rect -4710 2920 -4690 2940
rect -3310 2795 -3290 2815
rect -7610 255 -7590 275
rect -7085 255 -7065 275
rect -6770 125 -6750 145
rect -6645 125 -6625 145
rect -7610 65 -7590 85
rect -7085 65 -7065 85
<< locali >>
rect -8830 2890 -8230 2930
rect -8830 155 -8790 2890
rect -8270 2680 -8230 2890
rect -8110 2720 -8070 2950
rect -7660 2910 -4755 2950
rect -4720 2940 -3325 2950
rect -4720 2920 -4710 2940
rect -4690 2920 -3325 2940
rect -4720 2910 -3325 2920
rect -7660 2680 -7620 2910
rect -4795 2890 -4755 2910
rect -8275 2640 -8230 2680
rect -7675 2640 -7620 2680
rect -3365 2825 -3325 2910
rect -3365 2815 -3280 2825
rect -3365 2795 -3310 2815
rect -3290 2795 -3280 2815
rect -3365 2785 -3280 2795
rect -3365 2755 -3325 2785
rect -7025 1930 -6970 1975
rect -3365 1585 -3355 2755
rect -3335 1585 -3325 2755
rect -3365 1575 -3325 1585
rect -3265 2755 -3225 2765
rect -3265 1585 -3255 2755
rect -3235 1585 -3225 2755
rect -3265 1575 -3225 1585
rect -7950 225 -7910 465
rect -7620 275 -7580 580
rect -7620 255 -7610 275
rect -7590 255 -7580 275
rect -7620 245 -7580 255
rect -7095 275 -7055 1330
rect -7095 255 -7085 275
rect -7065 255 -7055 275
rect -7095 245 -7055 255
rect -7950 185 -6720 225
rect -8830 145 -6740 155
rect -8830 125 -6770 145
rect -6750 125 -6740 145
rect -8830 115 -6740 125
rect -6655 150 -6465 155
rect -6390 150 -6380 155
rect -6655 145 -6380 150
rect -6655 125 -6645 145
rect -6625 125 -6380 145
rect -6655 115 -6380 125
rect -7620 85 -7580 95
rect -7620 65 -7610 85
rect -7590 65 -7580 85
rect -7620 55 -7580 65
rect -7095 85 -7055 95
rect -7095 65 -7085 85
rect -7065 65 -7055 85
rect -7095 55 -7055 65
<< viali >>
rect -3255 1585 -3235 2755
<< metal1 >>
rect -7100 1730 -6910 2830
rect -3410 2755 -3225 2765
rect -3410 1585 -3255 2755
rect -3235 1585 -3225 2755
rect -3410 1575 -3225 1585
rect -7200 390 -6620 1460
rect -3445 810 -3405 850
use bias_generator  bias_generator_0
timestamp 1697389219
transform 1 0 -7520 0 1 2690
box 550 -2635 4140 205
use folded_cascode_differential_amplifier  folded_cascode_differential_amplifier_0 ~/Documents/VLSI/mp3/layouts
timestamp 1697388805
transform 0 1 -7190 -1 0 2785
box -110 -1580 2410 170
<< labels >>
rlabel metal1 -3225 2165 -3225 2165 3 VP
rlabel metal1 -3405 830 -3405 830 3 VN
rlabel locali -3325 2930 -3325 2930 3 IB
rlabel locali -8090 2950 -8090 2950 1 VOUT
rlabel locali -7600 55 -7600 55 5 V2
rlabel locali -7075 55 -7075 55 5 V1
<< end >>
